`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
j1/6cnkvbBL8f3aLllPvlRDArQFK/8TpKRBgndMXcfc3UnOgU0jGhRkD/YOPPvBF
2tftMgrEk8MuGAPiz7Gy8IzuDwyjYYyDsCpPZo7I+KVbO6GGEt2CyeQfeTFhs5CC
scgCOCFaM2tTgRSIqn4KUrv93dTeT0E0wfHcYbjYMLY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19824)
hAypeM7TT9/qcF6c8xyAYNidh6lr84lVPtGUyoCC16wJKljmJ6eVpDBxP4dnC6xG
Qpy74nf11EqvaGDA1UcomzmzK9oV4Hlkg5QEgdSuSL+FMlnCmVdcgNkDTP6kEvxH
oYcPTEAh7AsFByUcpEWUDTYtzcWIV+nX7jS/1OuubU1xx40KLOnvfYIeBBNhghzC
rlaY2BI1PDhfIuYd26BTtpllV4QsbW51dix1kGJ3Jk2OFfE//Wf/m2IacFJCB06u
+0uZgzE45VGzPVCzrDwo2is08pXCmraB92OIfclKYKDUMYOAylIi/F8xLRYE2cQa
6kxaNtr71LDjz59akSOthhhAy02rGL0etNAylSFNaeFsGWROAGoxK8jKPdoCjZnq
biQ8pbB/b8tDbxnMnoWELaDNpdct8nMeubcKaO+kKTRkVjItukEANUHh0WpNHPzo
BLoSHHwHLKDWT8qZvw651JTw30DBaztqGD4SyhOCfXw84w9dKhjovBO6zpR0I7YH
usNYvhHqgIe1VwERw/Pvf6vtW7oGzkNdrSJmt8DdWd2urRQr//SaPerGccUXkt5K
VOgUg0T4sPJZ0CB7os9fmhPVJeKIKi2UAMt+Q7nE5GE9K3iGsQXnUzZmNTVTzJRR
HZyQVZQ0/c3Aum/040DR5/PY/n8q69Kg/xAb1/dYiRWJqCgZtWA3t9bA7LYldqgO
DkrpDxtItZ3aH1jGkIWZOgjGbuZUzEH9/B6jCIcWOZxVPWqVv/07atsTgOyyrElp
c7Zpb4gvXcgfJff8t3uIlRbCNU7BZUl3vY79+29QkMxllDvrryP5feGsSQQNPpR+
R80wps5IdH6l3YL+DBCrYGeoqAGsy0qMj/KaXmGvr/4C9GqtZ+L8AoXJrx6leYwH
Q6p1n4VImvilzN5aKnHRKJhH/qHmGKE+lJKBiQv/GlpRvNViqduBLpUuPmycoO/+
KjgBRGTuhAARfKS9BbU5jFB0aO84LvQ6SY51PQhWAkgO3TazI4nWXCLo4FypdDu4
R/eZEwo6stn3m4b56ChUIaqhxkkg4/npd3j4jFFRlLBXK4sMCNwRf1zQ4uus2fsr
4OGi6eLtoFU8WYFQZ1OwefgT9G0mn22nvhcyT/5Innar3AsQOtxFqySaHRsPo21y
SxFLVmaUkWB0BMaun5xMTrztxES361klxTbSHswBCqT5yv6wFTM3HymcmvzL4lX7
SucfjVKPzZUo1WLlxKxy285Zve3AyCBFRwiwBeUFl9X8UO8IEiByXYZVHFae1WJ9
veO72rnUaq0EDSqtXR+FSzaX1QYD5aE62yPUqX7JfcFGBAQ6+iEKX9yMhno7BwpO
Dsv7JY8T8AAbP8f4pgjPL1hCVRfu2/Vwxv888bfUxlICHpYk4CkGJ6NbsVbgE0bI
RzmhDYBpE0qQCp3vQCDrxuw5cfMXDLgjUcTCQq4LtLdhASwk/2pxLpoqHYmB+sKq
ESEFV9rDoDJZ8BXHdwUxH6618aoUYEPjygtWyNZyLLwB+34WDQq5Q3X16zicEM74
Yj4pWpdk84YcgEo3qefBBzWyVGz3Jmlbl9Air5c88hja3vSoME4ZtAMPz5kIOB3a
j3acYLndEQ8vOnO2YSePs3/n8xbQH8jCJenOLvefGfE7j0vTUV0DofuGGzhZo2ox
54ubWU4gtx48uJRatajN7+du/rDJ3OlSTeGlOYmV7w0seZgbhYIHWfJKDL+Hylh9
vAASLgrdce8q64vCcYvtgcVRpMMHD/ndGvIWcdxFk8mVPLxPjqsuQod1O/sEWOCp
C6J+O2S9PnZyndyAoCxFJ6mn2AMuT6O9qnJFpTvwdzVABVBcZfJeYOlxavuWsBxv
cplHMilRdDWuCWYmgm2SJ2bJptd9Ayyec00erYjNDEvGva7OVRFgaBMjxBGAymZA
nT/jLnx4Zz1D2Bsutjx4KaadK7qfKRhmAmfsbO6KKa3x7o9fVubINfE2GCa+F9hp
rYj7ZLZLZKSqHOcfxsxxBJogb8Au7GBGYlnlfsCuz26FFK1OqTE4ZaK754BDrTVk
vev4tLq1Iqfncm5+U18ALgyz4kLb7sQxbN+GI2bGOY+t0MxyVeqy/lszb2h+AI/X
fcsmpNAgu68Lp7/Fec3b1GXVfWhCUu89VLuBRGkLkwidSfouhEGUePX+piDFitpV
1KuYORjMP6+pyIwkFfv/q677dFOVz9FMj993LbCzMW8yr4kkpqakQtfsmM3gom8B
1Y46Q7ZIGeafXAfdylhPIE7Z1YtPR2QsEaU7RCX5cMbTIjU6mSkK7WnO0hiJ2i7N
XiC9Xf3hed6LuSlsyW9dairKPx122/84fsMnxBqu0WW0dDolFE0yueKI9vjsWuNy
zD8CUZnsr0OZuI/Z0fkRydwYubCABKvg+n5ht6/FTtuPKKQuUiPbK0vd3BgrLCTy
KzdOB2moswNwC/mQs0eVvbgqyzapx0ls731skpIRl7bL4g+hvurm30dz3K6zpwpR
lIZ3hNyiuMqUrgHtDvslZmAqjNKLPdHs1TiOWZwdWbXhQOxRKlXWxCsmEQESzaqT
HZUWojbE7/i3DpnpTArn8nrDk5i85oOZfdfOPKA51vG92bRUvV2k1aLo25BHsvu5
qPfe736GgX0nOC1gpBouV94Qd6Bd1yFc4sxMRlgOOY3v3Ey9zyc2mN4ZbdRjiwNG
od7LvJXP0xzgm5fzNN8icTtGxu4kH1ili4VIAfpBwHH5A6MqGuLC0EA245F7IZ7m
pV1qiXEpi3uyfU7KEd1ebcUtxB2/EfHrb8BZi6ev3T2gykAqlZQuhil0PfMyIszK
z8Mi4PSq+dYlPAjxq+F0UHQKkrgjKl9b8G21SOR4od6zR90SwM9L/30NpmF6OA9j
ksyXcJP3zW5Wn32cKBg4El0P5oVI1Plyh3wDj/u+yp5uH9CjkpHhZdz6GZ+jbhsT
5XRpJXJciL+6hijxRfCjk3SKYk+tyG02+KJFF4CA946CbfFQL2JV1XlSqBtuQgCL
1IUotgK/MKM1Miu9LYS2CCpzfvF/fXuxte5pGt8i+O4UVexIO/461DBZoyqGuNfp
VmpNUj3DS14jTXQIoiNf71GkuKPvAFuUCum1UGfFj2NDjNY4LkyN769X0y/dgJO1
mCTu694r1Q2uJRlqkz5T3INHBGa41CIzBlGi6YfyUDS9Pln7kLWwcRvFa8qYA2Pq
NS1DriNkxhBXLoOb+YAOAJ2Iy/BDby5RuuO74CbYnK/iaz22d2uwZ3j+8tzhET1+
yOC7xc0PkK5zBlfyC4/heMdBUSQhZDd32mEEppJ8Jl49vUmOAMpeaLBky7XdiFDW
Krio5IC83SWeG6QdKgG6UTazVcxb4pBW1RWE0330Ex6f3nfONs1MJAdLgumx1lTj
uM6pFvC5marglQ8B7ltDrpwS1eaozHNdi8ALTYQM5QbXbFVT7O7lbvaBQkZZq1z7
UAZM1r68+piIbSigZgPjd+VmXZpA7hEZoj5A++YClizvRTRqX3UvMHWOjx6z43ds
hFqblPFuo5ve8iWgYng99ZyfuDvKL/U4TzHRSHO6thc8G6tskf7K5j55XUXDmihY
44IpR931YA2RwRQBQ5S/zM+NWnBFKrqKVYNTb8LorFoCeWJL+3kC+sjiaG8UvcJ0
BDQdd7DWSyMafEKyTndGSskaG2Vx9AQRVFjB1RZ5ft4sqqaFUC4aysQ3CE3+c6YR
pVoFoHc+B7d8zk+3u9DGPcyr5LdAzhVGaYQFxMC1wFgSBoWTi7m9GQrO89Eobw9Q
uSCP51/GfWDUg6HZTSsYAPqTzOiF0NOhMXyEyASmDm53ZvGx0hKF0yy9k+XlrLjT
g8cNjz1aFCKjlgGqK9v1WZiQ45Ujgvj0Fef5rhmEeZSw2tQnBqFnUqcYye6XoDjn
z4R5YZVaViSHhuZgxxPlc2jrMeafrKGJyc00Rmurh0tQwhH5+SDH+CiiHhxlWVCB
OuhFeFeNlAXoBntzeNFReai9IYGKPVnnM2VnpAlyOapnQbrl1wjN+enl4kpKqTKN
azGIgc3yQUGCYse5cP9BrxT2G10tzbjbrinZy+bXny4lXV55jFwM+7kXF0lhIvqB
L4sszIv/+F7IBOMmyL/iqRq/X+fGb4XPjILbW/GLIPFdAQdFFW8lnTXOmezjgf2O
pEN/tlymr1n084QU/wtvBv88SCScQzfqeF+GIVNWaZCkwmV5aQzyMaFRxSUtfNC9
tXykxnPwMcctDmU0r/jLSDB094Y+8WIb1/2ebmMZnBi4yXGOQds4ggXa1ctGahbD
1feC/wFrds2hsg6sPNkUA1KPMbAhQAvLeQSK/SWrGKdOsbfFXKPRHv7i2YvJInaG
81LYAzIhCBl/cEyOP1TBO71JSnI80dueWl5X5X16GMz0zFoJSLJiq+5TwgSXGzZO
7wRfz6dFR3YE8mgKzRipgJhCBlizKasZEPnHGXMrRQg8c6PoSF8sIfM6dKHQu0b7
uR1LSLbNDtuHx1QSkDoWOFdaJuBJlZHJSNmpUBIa8gkZbuHWvOYfvXQg6w+Okd/K
wKHFkztEufyl8eqDQIQ2fjeLNrSXomwIuEI/l4s9V5pFvv7Uo2f+TAN+k2DzrSbg
Ozdbbe9A5SqJkFR3/AtPJpUqTkdryy/rBEntGL5D3eMRExHoHGS8bL28MtVGCEuf
lDAnqeFHIEjAF6QXLuTK0tcFJjHU2G3/lo3KxFBk4uPpSEgbo3Gn2x7CI6kefwUD
3wVWV7SN7J1HPPI/ShwG2MH/37n6co3NIu+YYZSR30PNDsqBHI38pfGCuoTBE7Co
FS0VndUHZcCJbc4bGd9bVIvHSQBgQMd81RVoijyo2Pw9fae+Sh8dtjs//7Posxt/
M5E+ZhD+9xh0ddKK1V5yLPiKKrJZZkGjqt9FhfFQUjLnUzLFNWJso5n2mSxIE/gm
3ybDRyiy6ViJCSpE3fHOLukYM21zCX2hZ1St1pnoT0DVNQOih6Au439H8mpxc6QW
vVGWeKxKq3xk7HxKvo52ybv4b10uZQSmdqetlOC1NtaEnhLiQyXp53LyOzVcQtB/
MM9TAhJbMnxmBwK0x2Cozeq0YjoFmPQgJrhlq86J5ogHM86mFpRmYvJJ6nhNrhGj
gAvxledEs9ZASaIMVeNqHV71MO3AelIPVJBFcTNHPby+Csj0mIssyuQhAOQ+ej8u
W8M6hdrZiXCT7yeQvs4rlJtSoKgS1OhoXGluZoqC+4qslgBv0GeUBb7fS9tV1YdO
a0wPPnhIyOduYZT3PeR/pfs6NDlpDMdydZ8uMnDWO8fq7uAaGd1WlYI1G/of1SIC
Vl/0QH6QNRQ6rRBusnfG4qn/BpfO52zTCvWavCPVJ/fc/nzx65DfyP/YA7IRtVtM
+88H0Luf9+gA8kSoPLfGI1yIUUUImZPyDfUd/AcjhjFXBX9h33ESvrqX5nfocnZm
ihWZzrVhE8YEekLQzkxrChsB74E/fvo1x1WunCDV3M2tgyWm31jWIslxhtP9uNpN
ZkM3kwGUUPYWBfD7zWlKnz5oR/UvW3WdJwcMnACCg1sWSYHOogKZxUn5eroY+qOk
0iIuPUv9CJ478WXkqp87SJmLMlZVvKpdm8bG+2nnPJS972VR8KI66iIgYvODLBhA
eQTX5+WNNJyZXB7w6QCrIK1LmNWYG3TfiWhH/0g+ovfteBioh+gfpTED0nwt1nQk
JXFy81EV3XSocnBSyYPK/RpS9O2d7HTO1YgRXsdx63OL3FQDR6dQCOPyNKn5vs+d
YHjX+vVO0fAbfTOAdnLekr/VmSkBWJSWsgqZjw0xdkHdpQmPCx1tlaTPe3d3zQFL
1L6uyoFDk33+hjTvafy/I22XsVaupQI4rO6SqRk3v9SAB5nE/yqBZXQJN9pCgu+e
OuhZg5iox2wQHja2UMK2ncNBhUtPjZ0970yIH6hMRsaJFQDhtxz0Uz54t+YBGdpq
qlhw9uRtboEs+Pw8QnIKWnC0E/4sf5+nM/en8aDFIBxrrimk9P65KLWQmvDpK1Qd
yYtnhOP8WMY8GbLoX/HdIp33/P4qiSKU83lr1Fihisdw8u0Tqu3wO4mFqnuN0yKk
lUY+r4qc3BxdDt4JGXH1LZiOkvHNtUPPmxbnKfNsgaSN9TWNGgNnxUzYybvGcO+i
jCU9DVn/a7dlNSE3HL6vclbm6u2oTbUC58UlHhn5z9J0L1QUBZFjcWXGlYLasoa+
suYhwCubyRizZNWwIytANKPgq3faj1YvqZTNW/5M8DkJFqKQNjjI5LLZle3Vv92Y
rDt15ImY4TnelpyanEOcBF7xr7A/+uJUcecjHJoWYyGY3T00ne+LDZY7Piqqc5K2
/QdRMRO5JC74KzKerP8c5LT4WaewqwvvSJAnZ06gaxyrWSHMte7rHzvpDZxgujbl
Ji5SbrdKpcIvX7Uv4+iDvXBpJadbHD5cwFiI6o0y4/hM499wQeOCdObXl21DwJW9
FPEBdLM+YPvCoxbFIUS3gdPW2KzJ3mPfWqMBAigEAxvPQR1Ff1bQanE7vULv5qR/
XG434qo+I8E0Wrye3rTyfqww6bhgnBVRV14tnPM4+YF573v3WY3xwZFPB1nLORCI
cL8GnyXpsN7OW+1H7eiypDyMWzcijg32458DjBBqORvC/gQM/0ArzNpJAOP2JyVi
68rAQ9PvoVUuF3N2qi4ATiUBSql7i1nF3in1A6VnkUs+khCpwc484afhliJ7qpKd
sgkVm9DyEh7+VjZ/LosUZeXWkE1qQQzTMH53UM7CX0uOSTsqi+ZbYXAiHWLvhOk7
ieJL0QPNgVwvNLP2FiHVwZ6LHZCtRk0BaLE9dLHhr0pmhZfHPjYk/UAPXbMkJ7nC
aFH6CujjHFg5hgRBHpA9TdhL/CY1Lc0YvyQhU9PrH/tzYkRvUuaLsoYfQIvYu7Hf
o4MBFyc5S4yhG/ZUV+5JQWuPmj716LAcJ1DwLyhMoIc3b5Dyam8J0z1sn9H+GPbz
I9Jxn5s5ePE89InubPu29LSMlTMZ7P3wc39N4ipC2Jl5LhWU13o9cWQwMYvZGSpW
KE85ngBXcROHYVPyF3p7qqwgl4pMoo7yI9MIZ6eysLHRzF86swx9Hiy0m+F53KjZ
v5Sw9c2tSIrp3tFwzu6w3UVt2D2LLtfELxTYncfJKmbs8tYmR5bCfy1yadXTvKC1
u3wROxx9n4zF5FXjRIP7Mzr5EQCeR5jnDW0kvXt34tRvkvWycad5aVWwti4+yz2d
/MU8DM8OyS7U1VFQ4hhkGzMDEDEuS4SuZn1JAlTMknJuJm+iN6ncofXzHs1waXIt
a81k5CabYAnUdoDNtXyJmgCJ3zIeHWQLK0YXCjHN6vtkuQfzD5rUi8hBgehHNMGH
sptR9uNBv2oP6wltgQQFlBsLsjKjQOpcMdhZ2EGMHroCpzKJW6t8YUthQP6VabDU
+vSRSPD64HT0PKh9OIgVWufEIbgmflOFoSq9Y95KYejV8WAJneixFpxlff7/q8IQ
eGXzRWGtNbjZ2Gr38bPFgTcUWrsaXMqL8OmI+7cL1+idgSq9AgO0AkxLBXHe0MJy
2OcKeqAaVwXWROD+iq4gPjjwrpWBUfWBPNLkRvEtv8dNjUYidIJ1jbCpzrhgJGrT
eZ+m0vWRkEwbHogg+7RcfanMSyApKmzT7A3Z4DVoBTqx7ZBJPwIfzGioldc9n71t
cO8qSVx3RTmunT6QqMaz16Of5Y9tQNoSGtkUVoblcGEesZXj3FnUECwu+/Q5S0Tr
5Gim05t6+poRtREFNyMHzScp9Aw82MomyBXpEQdBmQc+Vx8G1vP9qMrmpdKRgDZd
OZmmzQjJSvyo7xC19mffhUmLpe+If/TBiCiOCdRAlMy3306qI556wjRrVt0NoUyX
mjqdWpy5C2lprcPl3HiBW3RWBq4bFgZ/6WNpKsw++D2Su2NNTTNToG96A1XGpAJ+
mGfWhFzrKMgWcpmXHUOEHosFd8pnQc7GYdFyjW+LSwYjALdUhDIkVbIJ/RM1l9aD
QPXdAkTeQBRFCJCx+v1I8EMlxGWrRAg8akTHEeko1gp1bmzZu+m53Lqj5rw8qhB9
ufJN6spsOXqtTpryRqc1BFyDZZR6KNTjTmY/nr8j8LWDke8bUoAD6NPiUo54HDOj
qPCcM/3UUE+RBUEPu91r54fXBv4asdOw6QTLl34RIlU3VSaif1qmbrG8gVHrA/2R
AnFuLxqyiOtvSzBhDD7XIVLB/VVMyJRrHWwgAVCKsFMzRURZaYGInSCD53qQtull
xoEf+k4e16gJxBhoWFkaFUaGCbuRqk1dUPzYMOH9yEONqqNDS+H9/d1zBHn/X3lx
oIPSSr7MWHQHt3rBC9Ug/AQ2u3/Eub1JASaicF4EzQWkdqBFQPEr9sPMNLftUSk9
6PCsG8DioBdD1E0vHnxuCQCXRrZFlp8Q0WLp4qD0oPbD2PSQcGtpv/UYTnnTi9r5
V55wnnEN5tt6djoSHxAUZWa4qXlvNbiYOqiiBtj816rg/mauJliLyCELuec6zI98
+uVt0Fn7ZNRtBJW9dOgaW7TyN+kv8ub17zwnLl432tuAzz78Qqqu/Wv/y7n4RXwZ
QBqOPMJDW/KNU0t6A10d3NwtE7xB/bi5CsgXdlz0Lzyj/BknC7ZYTqS+if222hwt
fTKCQrELJnV+tppFNkLAbOj8E0oLsvK/ZI6ChhxFvw3usuYfY64kDWvi/zeZfyUK
pV+JwDQIFY6/NLwWoF1v29VN0PAOBt8oRL7kgSR5ori1Lc3JWQ5blyYEqX1H0ikm
3zkBPNmBBqIcy6EIQFPOaDsC1msvpU/8lJSqh5MdJoV4+2SZ3+0i90Hvp1L3tixd
WR6dU1YhwMAPpp1u9lxdrcFWQzH5c4l2GBMAM61V9+cy63mXpxc0+s1cafIhHjAq
eKK/cZ9qWv+gtAejGJ2B63l3lLFGfehFd0wancVj552EjhF2uTWUPJP6YH95BBBC
aLldiYBqCVxOXnZzgurGEGSYzwvzJHuuiTPpxmQDhre1XEMUiS+uGTbTishkwwVs
c4GxZnBwK4BzApPHf1LDOJo82Dn7cNl0GVGKmt5ghJMnWhous96KlyoTkz8srfg/
KBQVr3/yiNvBWB1KctFzVdwafeTx6X2y8hsC+iWxPHUWgE3W5QX2Q48nN9P3YMOR
fft8n8ImJ54ecAHnMRxNHrQKaMSo+mvHi5EFgT64Hb+6e/M2Qq/rBzrImgYoWzjm
rfBcG0+EdTo8YL3vYZVxxMTQ235KhYn/tt49OSCS04GwO1CnPo8M00JHReel6+Mu
YrLNbH3pavrt09GbTBN51caF6hBkStYw2lgl0pVetpUMs2J5z9xhfmEsiVF2q7uV
Jo7piMGs4nNM9etp8+vXfA0Cgs4S5QYpqMCoqQ+Qj7p7pDrxjtNNV/0yJxE4H3Of
NPnF0cePqQ/xkCoecychD2oaDjx6bNv+kQ541ejKyR75JK+PbN8uWuzSIoifRwZ4
KLE4YoL6JtjQFFvZNCEurjlF1dnjZzEV3YEgpuAe04XnZzW6r2xCeU31Jafblt1X
Bq+N6TKCgAr5SYVVQyinElNpQk3WVi18mRLOdCzzvad4UO2SNvdDW+cP1J24sU/o
pVgK8ovTuKkF6WVpfvbkNgX59oNiZNF/6WPhQCNgPHC45hA9ZaUehi6uo86bGESQ
Cr9F2yFosVKIPjF+g9x8tg3ZWiryKCA5cEzgmW79yCW4Hb7sQ9EaVF+bGromi2ZE
1WwSgrjTMgpdvMX8SILRhs4unWnULkWrCeC6CqAh5YcK5E2KrUnn2EcI4RxPr4H4
1895dHbsjaiqgw1yqDuP9LcsMcf+6T81502tbGo6cZ38lLDgPoLpsMdn/nzbnK+K
P80ACkUOIfcddaWZqLuE64brQLkj+Cro4QRKsa6KAtPVotFaVZj4nZx8BI7ABp0n
oIe0GKg+hyY7kEAzLOr2LyuiAKK5MoOVvnyCiERVZjdBvzs+9bL71xOmm+bVWcq+
57uH5RXX0hjk2eTN9oaWI/jB4Gf1JtZYG98Z+/+XnmZBK2GE/Yw9W07OcIMhw3Pg
wBnvRmYbt1dTQ760TslHC+1b6BiFnKb9kdXMbpOb9zhVd+iFHvrkBQKeCylEgoyd
TP5DxjpNBEIR2D+1r94vvrCxEiX67DgAZJKfvqZyjwuXUaYG6ZgPojBoH9Mp+XER
q3RTagfPuBjt1X+DxfnypUdRapzqPCRphaOzD/V9YvtuJEE0xHkY5a8GS9X6Xdyr
w1KroO5b9rr+IEN105Bov3Dpviu/ak4e3EcsslHiMN4amU7Av42+7X6D4HOuQrkA
TfCrAcTG6JtdqBZydBn7HmT7gBEC3AsHE02uFE8OrU9Qe42IzqaioG2mNmnMga3v
aI+9DGkUno4mDtvKWkgjvJibFc4v4LGf4STxC3xJJPgcE7KDgHMRs1OcrvOgLIKn
t9c9379aOYoOZstye0cYbrZHNXF8RZRVEcVcplPoI1Y3EzhCsMCZNIfaDBY4DOlF
HD4818bWhJuKVXECPpTPfj2HG+3FPirv3Ki2OLvGciEh2i9LBtmdUVsTFtnmVVWc
8PiHtiEDtYusFVyO2SQFSRJwsrlqIbOgRm+YANoPfQgsTiAo0Ne4pR8K74iZEwVe
rminJkqJ2Kt501tg6/F5U2e1KWTgTTkRqm8kZHXwa0apQS3o18g5yPxZjb4N/KJ/
L3WetPXw9rlA6ak0v7vNmAqEEuPxNzIiAiILT2fgK3WiWj+9d+Z4z8NrW5z1RF4W
Hi3+ZlC1ozjgxRFghbyOKhW0UJGbjNZ9c1FD2VQwCKwmzs2WWf3CE2JtlgqfSnYx
Ee5ClGsXx7PZ7pGO31lBElJDTF/+ga7FnPSwrE3jke7Tvxfi/f8SuvdZu/hOs33l
HmErwaDJfWYvSmf+sTzDAWXijSLy+SHGLLFtZK9qZJGhi330/BE0c5w52QpRpEau
TcoY55iss/cEDqF4Vsbqnc6S/FZuZx4/wrzWdTCB48+WV1d+VNcAlKHpNx/d+G8X
0udJay0wm2biEHMrjSIHVverFdFa0T4nm30YU5ecov0D7Det2kPHbM+bDUfKV5D7
HUsvifyQh95HabIIo3uLFaz/xWJw+6rWhAiG9agL5aq581xpo9Jymc9mq6Eh1nw2
pTissm66FtRyUtYtH1kqQAD+v4BT22CFBZx6RDxnCihY57CkBX/NHvuE/vxvvuJt
TM+kfJyBxVZ5TGsaB9Akt5yFyDgFsKhgThB9qHOtbgcz0sFNeCGTWsPgsIl95b/Z
LwZUevQUlROUktAw6jFu18DuigaamNcGlHtMWhfgMu1iuAla7MSINEJK1nCMPau8
6fCRtX8Gh9EB3KiMZlsHpQXJP7munzSBmoHdfeuhd3x+UJq5BeH4UO4ZPlNRC/5J
ZlJbjPRy5izW5vTgTzi60N900sNQVkla/kKnNGCxvdiHeAWGFL7A52w5lQVZoisM
JbGCk3UI46m2U21SUsZrlO8q1HuhLprO6H1zHjxFclYF/ZIHtRfei1BXVf29ziGk
qKrU+GJ9wI49j7NSrfTC0W4nAlt3il20IHJVNct90+TkkEIVNJmptf5XPkEPvrh2
KeUlrKh89emOGDvDu/LiQMH9NtCOu8iNPGDugXzv0G5KwN8dg6HerGtKlhGnKCIS
FYlfJ5PbQwT8YMXB2rIcmnir1ibIjvVElTb/QL08CsJr5W2rBl8jRU0GESQeEOiJ
i7MzTOOpc5vZDoS5HX2EJ9MqL2IgLJ/TIIQlY/sGxuUN/UuziC5Z8OV+svxty1Me
N/uCzztulEfhPeqC9hFZMmiKL421pZXni6e+k7Jtl8E6sF3vLE7bFs8m94rHliKt
aE5aoX4BEFbJz+D2/aeFYLG/SjXo83St7Mu26r7TnaOXLIpq7IzB30MSXAIojiPz
DO1jUcDUAG0f9kSBbKAQoykOn0vUJThCX+REF047avycVulrk7ZVKNrM0bTWCZis
RCwZVWccVtAKNpUG6BKw9zHcPDz88eUEXTpaM/8fGlv0Uz7k389SJIGuSopJlYMS
Z0P9zh30KG4cK5e7g6hiFhbtJp3w7CWDMwNeJYXC7zZjsr+yFyyZFF6+Qxj7Ybi1
oRZM6t16DBxO8gGUDaHZnAaXx3UyefJ+zPrJXflp0wqM0kESSYFV+vXINca9aqMa
lv2vYVb8V60nxiywauEJ74tEYhWIfyQE5Tx3iQ8ee/hPdWsolHozXMdOeIm0AtGk
tgcoqUyj+vKeiQ9C9aMB65YhM7ATwqGiSVc9yC5sZpPPGlc+2vD4L11K3AD6i6z4
TPawfVaD/8TNGWCBlP6MXaRwwKLTJ7Hiu5vJJ2Wp5j9dTmbVdASyMx6KRD1GJ7PL
gTcrexzRmjbxYDXH1hYzUyeISAXIRAEaAcvGAtuAgy0aU00WNV97KBDNXefN4Oqv
1IKiHPq6ShjRf2qFZk2wNH+dB/31NFEEONpwWQomKvvthT7H38+bifx6jp2EhN65
HyOVwLVicEfGJ4bsljvTbOr6NqbdHn9qQMVDLub0EkvCuWp3VplpOtUl26v5gUpf
1yAoFM84p0XYeeABVYt/J2uXCwEZwpwDz8cC6IAlVsEr3mlL4DA1y7ciV9y2Q7Tl
LgngmtLx7dJ+NXMjpA7IdIsdGWmNeDmNEA6TGhxkOw9gqiOOfKVMG4n6XdQRdX+t
EE0IxXnY9mfPTvqLEhNz6H4c2L7OLH8utywWGyoaOz3S5YezsQlA0HIldlL7XnI5
ugvUP1m6qp4zn6pu4J43wtqIpgKx9VlWHP8a1aKOv2pkqzFs6CCBUc5uxPK4sX55
NfBWHTwE4pftQyf+bv2tixurswv8dsllnQVGMjOIckH6zbypanAqsu1UsYeLtX1g
n1du0vQRYLa50THHl1dyu5A2Fip5yzsmC5Nq8kVr+qpQsTYpqpK4DJazy/TtdEnN
+NXWuVGxuZimK4trcw3uwW5LC9YyU9ovBkSPHnjJ9gVY/7Q+lBhN1/g1HxLmM5EF
DvhSIxgSMYvylPYPWb+vZ0C6qS5hXXZ8AiTZmr5XQvyhxSLy6BCTsAE7YtxKoaPa
XV4xwBskux/FWzl75+NlKur8S1A9uhzzKDgzvOCs2SA5TRk3d+BlqpVZrqeMk0RC
tBNft2kvXQlLto/7BtIriXLEjXm27GlBZH7rG3e/sHVvO/cZqxNSSi48Xk0ru6rC
m5QJCUE/iWtgLA6O/TZEjMVC7LLqQw4DAqBaYufbwd6Z0fnfW44fNVXaFCPxI/gm
B+I1m6gm51he4iC+O6BoFridFzhxNok/IdWxYfmEtXpWrKaKv5dqVlzstFo97JHk
/k+4JQ0tzuY7BVYhK7iElN9Dhxv4VYiSd/UI24YWoIlXnMnGNjgNyWUtp0U+Wq75
LWi4HUkqdqyTJNvFV4emK8XGt2yO+Wjd9OtP3fwKwZDSIQzcq8j7TpQq2N0pF99c
ZNZ6lUzCU7dNvH2pIqytvQ5Uhj7PNwQx816kzQ489q5yYfbrgS0YUo50TKAyld2U
lQMbKOzbafSiOqbpHbk1e//jk/IkVSv3c692SJsvA6uRshYe5JcyjR8N1iZYhVSs
t7AUTCxtTIF2OWmKEaEXLOKlPT9I9VLENt+NZQqAh8QRTIqyhfics9gRbhE9o4xE
GUYkbLjgKUx6xRWwF9ndX1nLhojpWm8CjKH0gKBaFQ6JBItOidxqqFBV4hwsGo/6
pgKk1Hwq8qxLwluR3smsclG7F9r27ZZa3a77s7/N0nN7nhrjkMeaBP7HJr0JGWq/
u/i2y9b6SitWOG4ujr4ho1T1wHR97+eh+bBuaTk9bVjilNsnWO+zfptICjj732+K
m8Zlo+y8+/5oXFUAf0jF+EMGxJojmtd1V+Nozh09fOGyRNeA4nSMzgtvMb/azyop
5X2OH0cP/QUlbIGHYOI4/uO2JQo9IkFS9KrUhjY3HMt07tq3YvCp0lcfdav55ESx
jnz632U1rkZPLlwiDiNCpiV78oeedI7Tt8PlvUz/8ISIjVTrFyrK/pCmO/XdB2ev
MXT84aCmsp1e0790JXgUMN44qW40V+kri0dmpBk4C6PUORjNAYa+FzrR9JQTOF4I
6eua1lmB/wlAWvZg77oOjGaNWdRzpgH0OnZ5IiuI/JbE3fk2ydUZECpKmi6ygWem
GyrEUIS+RG6Z3OltckSssvuLzo9ZNV+El/U0rLIsiL7s3w4h4E+r+Tw5eIodzkGw
YnWWWh0c4uaQp7tuIDeDNTNvRs3rjHuBzQXyInJ52g3E5k3xttovLyySHB843PYE
gr4tszS1PpLpBtZwsSj9l+x+lAK118s7qxMCtFgQmZMWvWEX6HAe4hMTqr0nqbXc
zBjFO4YmNeiELHxZYHJ732oWPv+JWa4WFG9BGor+cWQosoudqzhq3KE0lOAs5s+y
QNaIJ901k7LA1C9Q/mHqn/65GD/0fXnq6ZDcDTgMWTc3Y6KxRtCjtRztE3pkdJEb
u9iPu+IdjOpFKMlXbQdMPnrVeBiqiN1tv9sBdnPbO5Rkd845f2eS5jf15iLlccW+
CprtkpsNQmxrIvnRwyrCKosLoytyC5Sn81bl9p94Ap88aoMN7IYR895gvrniGWwJ
5rLb1sb627lqBaUUg1YllULv4Zz36rhvX6Od4hMC/hdD7mNX/83MlFTBdXDSR37p
AWXWm0BW/a5K2gttBDEwYshSp0h5gzfjuOexlP6LT14vMBHQMvj+hrtQaQSjbgXp
vvWheNZWHKYFz3Vpf3qb0NAAEzc6eT/T2exrhGW89m0xZz6UnZBCoitAx208K+Vl
9sjSUSlYxqiHJfqjzzsm2qw2dmiByeIRXWKMGKgHX/TVuXJPLx524FmPuqmhUqUR
9Tu3jIiXqWC3nWt+tNjlFxf517sVe3BrqqI6jphIRGPxT1kzg9YOWmaHAQsO4zs1
BlPjG9HFuHEp+nZQK4zloS/O6EoJEaqTbspDteFL7BmN6R+HCWxBpj87/buWpF3r
+5RpG7cPqBy+ALjCG/9XRHNUpyZi1/tITEjBiyENMNJeUvUK9wpq4c2BqomX7IoH
EBq3doN2VMYkDiGgi7DVBNW0vZy63lyAp4zu2HhNN0zlqKKZRcRVTLsX68UzLeid
D0di4150f15cMFWzQFwHCFUxKpZ0XHl5TvGT8Hj69YiC2BAkWa5GEeOukVrHwct6
Qbr3ak8kFqW5o9kLTeGKf+j9vhbMUYg9CcciE+cxVZJfe0k6At2i4/C+O2ewYGhM
Gu8UQ/XeTlCJnS40pU7jNVnQWqmpzq2MLjCH+yDJJmR6SQXKVtyKshbFeuRxo8jo
Oeg2JZE7DaTRlgA4ohqniloJjEJR0skTRTyu0C3o8RkOKADj0iYy00xU19LfE2in
Wqy14akUAA2Dt/Gs5K2CmuhTrGWm8+tgrF83gt5VVLqP8RTwUo6HyKHzOwr/Mx5W
YgYGO2grmOi2oe+8mxocWcWZ/NycUWuNpEtoS7YcJ7P4I9maIEyZknZMeFX7Djq8
FgG7ACTk65dEDv2IECJOkOLiXQXYmkfvo91VIYiLqja7SFfXwmkVT3r4wDCzEhxf
SXVLNpANg9YhIC/D2mFFpvWkSwUCkhU199RF7x0yqE8Dtn75eOHco3Ognk0Yyi00
CJn2+BaKewwiqhfEATBewiGKZoKwYKOqXuAmGPYAx6u4p3SK3a85KqG4k1Seg1lZ
lVeGVDDrkzEaLIWB5MgjSHmr7T2ANzE6EvxBt0ELX9kSbI+iJPPdLk39E30xCleB
ggPzi9El6LidtDCPEg/Q+gYSKdS0N3Kbvq5ZmQuMm3e7cya6RgouU89EEtWBoVgQ
dqTC+k/aRRxEiD1nvpzP8HRzd9374+hON4Mx2U+0MplzLAgw1E5wPvyJdEFqyYeB
GWqmqo4sATQhCWvVYMeQ4L5FoEs2uHIf8fdu9v52vDkC/YiiUIZrFaRB6IMKaPYE
6smBzhIsCvJtUHH44u3ji/5+fWGrFoJEef+nFn5GgviPd4ag2h+7X4majIQn1M4T
EZVQ7yPh37z2uIQD0hBhT1KNurSJgXeBty3tnkPNDs6aqstOd6IR5wTa7U3jyRAX
wUVd0ldMCwXulid/jootctXiW5YZmgq+6/lomp0g8pzZ6B8nzCOQz9Os/+1pQYrN
jN9/R6aAiuczy0MZjGUFHxid7IS9zzkHrCyt+aY11eYGpCzZmFH89exS64eJX30v
vyhVIJemjeOQfiLRG6iS9a8tXG+r7k6uOj6zb3ZQAddA2BLEgmUCAMa/XQl01O4s
CIpv6ZW2V8SnARIaIRWTQMPTBoVpWuXkLqesUGiKYlogNHR+3EAfK/VfEYtkqbKA
3fMOdOuMRYQdIULWYS1GcEWTjcQg24x5e8GKRS486ODtLguIErJE830Yf3KJnpzz
lUvVeUmJQQqkcLiNYHttNvJ5wkX6yAc8tNHx2nZK5NRJTmeUMLiRZADBpaWpy+TC
7ngf8vYGPOFYElMixHiagOrPXo5jPrf3UvyXhvB09R59GjepbSjvVnuB5Iu/9cQ9
3BRoFvuiHulkyKqVWNwtoPEvpQkhpaIJCyqy3TmwVLl3PPn6Ctuo9bFilhbEXFh0
tTN+7tcM4zfk6hpuRuPkrrSWeSu4uRp6uc+YCP5KmpEHG33fKJzi4oNI2vGeiu0P
zcP82XIkYueznTEvh7z2WeuT62p3v/PdL9oD3ESFYWDU26vH44NWeKsSP7+qpySS
Z/OyHtPu/X4lK4O6J2LQ8AWU4t9KoP9yPyshBetW5igF4hPZrLWNZULUskp9yMYN
Dny54Bmfb8aZEuDATxGC5OsDndMx15dQA61luiWIerMCjTMPstryF0gEWO67/zWb
F49sP3eUmYw5H86mQBR31nH8v4BLrzw8xCd9oWSoShGPAV5Nph48UbqQZ7qSKGFc
KpxBToPrheA0AvX+WaHLH0sYD5L2HMR2xZ687qnCcVLCK/oCZkeL8Kn43UyZc1QN
y0uqAMVxvF6Z2sRX4b7cxAcRTdym/3TYJypDBanpNv0UcnG6+Ot+7aJJEXlJRtWl
MhzUOKRxRnfFdxU85WN6VfZkn78EgEp+ihnRnVNva+Tcze5a0eE41dQmOXhmvLYJ
XU/sIwfoVoPi6d4106lx2PyjtxQo4GDeK9DIvfgsLzO3/1kSiUDLH7sSD0FwigWM
XCO7PbNlD+3Yb97rOxOYtc55kTmMBgvHqQOcRBHGQ18tyMIYofzMyk1SAHPxWQJS
uW/1dd9M5APpTQGNTOZUh3ntQ5xfFmWv8mvGBj7VEOqOqlaYv577KDwgBfrV7wGn
l9fb9cl1lQst12D7pLqgtqx/avWJMKm4ASzjbFCBGZTAVa/yGXKzI6soQX1M/Tv6
bXvj5FRcGq9gyxgig04N4rYFV7gz7V3lYWJt0DKBnGTWYZgufef7I4fiONvLfc84
dNtuDCdiOOQ1pIcCMNYTDUSrAc4/WN8fHdR50CXKtHsgxiG/fOM4g9EPOeXLK0YP
rSv/Rzc9hTiI0u1cRAdnsQBwCmWH33e4RV+Wae+mzHpg5VLTZZmHXFOIfbAO0zHx
iDX549PZldh6pWRT0qwgNjq0zuPKzFG+JUWlCX6e+g+20b+RtZ7LnALKuQ49tKlo
MV3FJAA9s45Sl3JoLtzWg8sJi0W9pAYFRC6xN65sF0bu8FAoSLohoxR//cV945xe
H6qxMJXmPpsu5Xgf4tPuN67WMTlqIZNZGa07kUscf778qgonzhVdFG09iR/O6i5t
+ViQNjl5iEbyu06KfkFPrcYd+JEioflKNswM8B8WMb/BkMMzVIcC6lCzq+/1jjmA
enmg0H/4iYroU5JBjDkqxCaXSQc/3DleAYvQpTtGSmgCk2yQp5BbpV74NWcxsTWc
MUC55vgaCQmOMFwKBnBOhhVc3LrUNF9LmMQNYa3pAR8n2GN1VRUFrIBBxFW2u7Sy
9XA3/oGQ9XJ+ykghvPxcX2F8hIqqUumzDHQE8iBnpFHXPhkWPmDxFnWCwYJ/uujf
tKSD8++kdubIS52u1MFPgughC50NYFCDxhiWvrCQrlQ2pFcglh1qbwuVoZmq6Kuf
0fPM2bevEy9VIPlaOzs+svgiBrHkxD+qBAL62tJZd0tHSTFGwPEfLLRDKTuXjWHI
+cuBN2DqL3VpPbu58b17NuI3P1npYfhYOKkl/9mSlrs2of90/u02yrxwhx0hfE6i
+F2p9hVOa1UTCRrm/cN3zTnD9CW5ZLcS0FsS1s1TV/JrTWdG5Cc4n9JfS2nesiod
Je85Z4jBpXd6FetSQZwXUHe0I2i1xKIJGEwUkz+1Atq+hGur9EQ9QBGAyujAz2XH
HrxBVARafstk2tDGvgveRVumrmR6iBi7YB1EMcg4zSVHIOC9oP65x0X6Y7ULWcZD
W/0hETig+Ro4phFI+qeJQJOUf9EGkVhfUk2jd50jgVr2XINR3vZ1oVkEYpL5gQkT
4wTvpvPI34PWq/6lCT5Yf4HIcP6vc+VuCDRBPnTok8ak1bhefC/DqbTzHBqu/2m1
yN84zMrcPr1R2MhyKxbq8dNwfbtIgEm5XcapQ+7k3A/fU7xn2MLNlfe0P8dPjo7q
diDsRNDdgDsnQulPLCjPq3Wyfjby/2SOn+PBYbCLptxQforAr1yE+jgfJ7weJNnK
q5Oi8WnzlTSTarQ1yzOR7JdXntXjae2sLywSgj7YuXQwlfKblXRYEjQTFNZsa+EH
tUihi7NB99nGgBAzrIxYKjjJqEsQNbmT+DrMtVHITxK24xZXOnkebjc82IufxGJN
aquHLFBLrTfux3o52v21y/DmLqGNJdISCe01qOvU+ktC++vLW0bRuksuu7M4K0uF
z2E5d05dqAn40gt/j/Z9Rgug5Bd6GfF9C5Z85af9xVJiE2+idi9u3sarmQ9Q4h64
HwP585r9lM7UKTQsOHkETKi8KkTZZ6BqhwN4i0R3SSuOTCA2qiNdC5sqdclfyphS
7UWbT8tigDWwrR8cDmkmVK6/w714M4TRdWR2eeachsiXIeeA8RJZ7jmY+ki/oXxQ
TQa0G8yh1xntmRwWs0UnhjXLksJEunj/1HSEmSddS4kMl5Jgyr0THvg7Doyl6Iwi
jRA7X7e16H+gx5hcYidpF9RURGaUy1uLnD7hmCVT1ESAYzJq9HQqR6PCGhGxHwDU
W0CGxVx7FuyT1UiUnhvdq6F8uUYFNDji0ZaJ2siT6e99BvVwgvApGEo2kgftKOds
eVzbLaX6qPsXBMXP/qwdyVDZiMEziQmUEYG5HbTx7KVvJjhurxckct63YUgEL36P
qHuHCBbVE+mHuHt4CRwmfQMn/ecNTEhmMiAZcIAriX0TLGzl7MBYbOs4txYI+Wcf
tGiLXLblPbMMHUFep3/w+WqQXKXI/urK0xLbiBBTeTt4JWXJ3BSoEOtJ/Ab35AMI
oxpua+Uf9SM6spQuh0L/W1/GbH1UsgjOroewPMvwYbrBqtXw3FrYaMp9Eq4xEVUo
5rB6jnHhl/jlPIii6iU2DPzIsmJAe3ZyqemYQSdokcRne8JPKhwiO6NLhWqq6VSk
JiLfqeKoInGFDdctOsvyHXn4J/fy0IRtz1+PgLsuM/HaNxNopROKgVRZgnTGMNol
qOkREp5UoU/bjugfJe2DexcnnYOJU9R1R0BfEspMLJBqJZ5hVcL9lyUZliJtFQgr
QjpC0zWwzmQdEJfBoSsnGGutf1e0syxDdNSaTWnpevKQT5bcTZMqsYI/5jCrkg0J
Ad6l10bdVutvzwoJG7PNoc/d80RBeipsXOqOCA//OyQPOhlmWoJ0KNbvW7zYcQvW
qWLQ3HfznN8feUqrpauKGdEWtdkBH4C5Iqtvcf0jbc0ZiiU7jxwDFn00f/r+7g6l
kxGcZygfBJmOXwrikmLIfQYecPSImRMFEcqgqW8KswiPZJAXyBHTZqqPCw/hmZpN
TzYv72AFSDDVe88GVO0wA40RpU/ggsApHicJ4yIM5nN0bQuzPSeW4X+b6fDqLulC
nXhXT1hb12J288Bf4pP/i0ScvZsLFIXR5P8xbQi95EJDUBEe0ibmHC00eKLZt/AG
VXo0UiT7IMMSIDSlEP8vScrPy8Ryuz6+1bN3V4nwC3nfGx033DlUWvxr2JP+Mx2J
7IPPdzpbOA8lMC4Al7zxtUReVBJBvgpGk7COH81nTx1ClFSW/XishaNKCCctqj78
HJfoMMWIC7g/h+CDIcecyyLVZBlNY8JKy6doHCzmJ0LERF23+bSU3eP3ECiPjP37
wIn+2b00j0YAq3tUNUFPHo1bgbQtLd15UHsJ6ekKFdBxjgg7sfx4ug++f6MedJRZ
cqlQOm0XRXcy9mBR7IIdsVZFKlENXA7iwJ3j8PLh6YaNYIK2BBaNIY0uOKl86BMo
Eo9mzCjjyzqETy4tbB8zNNljI+PTWxhHJTH50ixYFUle4xezZDKl4LOFw2mvUl/I
AXGRTv/ySrkrISa3J238nNXkB6RHfQGbjRtJqDDLhIVZP5HcSONtMAmeWW9I4xmD
xK3ffIPIvDko//yJ8ZvvhQ9SCLRQ4XkCBsNHltT48rare+tf3CrZUXIgHYe5Vb5e
0cZBitbMpVMZCZx3kYWxa+/1OXHgDeWVCA4W4/+/+osEuiFr9x8HWF8IGIZfQirh
n6cAMhravhEAZXmEvNgM5W4WO8jWFXAUAuaD7NDNlT4tBIjGbhgGExNqjSBwWgZF
xmgX2iWIpJealk1UKtgN0NdEE22jPWKloR6Y/shLpu+sdModIyEsBVFgnCkZp7V1
dAKa1orImO2NmndtL04pWqv5J3e78ylV8xLVFcwyBMVnxv8eMkOhBvYNt4V/Na/Y
8EQN8ZYhpqvQunOKg1ZglxGoztaN/N8Nf3FrJg8K4s/IL1HNWgRSk6eWlBHOBtj2
y2evI+qQzyKyTqDYzQkwpolVz8bb6FP+qYyMt0wMVJFiZE/eWQVYb9y0zVBPDcgX
gcV6XyYM3qY/oHWKJ2rVoopEgvDu1H36kizJeVpjYU88vN/B1sKltUeFra0GkHC1
2GxyOgyGOk+s7qnj29jacJACLCd6Aq1emyA58DaaGTPN972uHzfbvmRcUi+KLgLx
jSa3WsDWgO7x3DktK89UTb/EgDbPMPU36BFpxL1akTSvEH3bEwdu/JIiDlBT242O
mL1/gwZCeI06vdN1LsEONkAkYm+X9jku8gwUEBtJqYT6mGar3R4TfyLVSqD/zg1x
TEbe6T1gRUt5uUBE595hQ8ssWOJXd4bciwUj4isbQoMIhYz/ir6/8su+o5STcSUA
VDbSYKca4fOAPvaa5bStEttu0iRdbf/k3WnzXyNjFwUqzCZzeKXXOgBQXn6HpLcW
lJl4gWPSgfHAbK8YMMlB1wfodafr+OcIHQ7qAimGBa9pPbbQhN+c7IxLB4ALQttH
9zwvneoaHLEY2wXCneLo343vbSBB4ZSODwfHEoRi5mP15QtcCL/lMfkJhQus80KT
39CK+lZt8vozsRXCFSni5e0ZherfuK3ARDB0MxKotGsYTwSOusBtfV6lGW5XXTbJ
tEkFR7PPAkGCczNV/wh0YVD7iWUYkWAtrdNpFL4tosNvQ6w3spzovt6VynCOW/EY
3WyIDUeAbBI7ELXdT6UfiVF8dkcp2Q2cQ5PFRCpZ428NqEMf1XpnL2AWzTPl1Dxb
H4C8m7dUzKX8374ElxAX+f7Dml0yZZTWC4JcKbkt5NKbcEwlWonEBv6mMOGCXaeY
LAaBPcxH4+AMgAmXhjLJyyXDeSlBP6bS65YIUnGbWzTpCwahJFaq+ZqTfzGO3jCT
2SSyjVqgvCdlFKrjzp/t85w48cUr4iCkAgnL9zHMaBfkrzHwouItnAZPbX/zndnt
d8gA35YhQZFcbsR8Wh1hMoMf8s3ravFMQKXqea2e43qaNNoPYSUuQC+aNPZq8/wA
m5EZO9bvevDdyIy/JBfGncN7fF7FpsP0Ng4NW1Q25eTFK5zWBi/mUumdpdMqv+mT
llqna96EwEH+gn/BqnH7Oez05Nx8vBJMUQXAjEvOA5EtGUUqelb8KjXQksEzOXQr
wuMDF8VrIqDnMT3fLc1zyPZDdXBtDjTDcvs8zeHLkD7wiJPwdZJTa6qZqU97wkdC
j0I5fn20h6fYODhcxQe4ZrJN14HnrJu9QktHMh09v7pTZ9DmZTidWLSYvhbziwfS
YYnq4cWVPrOVwGfmgM2oxWw8ba3d3fb7INwTRzDS39vOu7CkjM5H96UtpjCMayqA
BnMVs/jntCmBTtLX2onq427EBlCbSK5rlQKdkE8krmZ3TrlETVyLzqE75iHo7NER
YelkZLgiBLWQvNNyeOD1M6kjcgsgbFvkjt92ZhBlzu4QrU2H7TgAgWZik1B/RlO/
/oOQuIXRSsYdu0uUJgwWgx276VS/4HKoMgqNKgIeXheGSbvcamwtKqwqxAB6fs5X
uMRrR5vm+goyAMBWVt4KgdUedPh4WZce48spmgYZQAdLPLlAlPFmI6wap8qX2Y06
FzYYIgxlph76m4sKXlHzjYb0jH/gSV0JnuFXjPQOzWyFk371mRZi3H+e8gd3VJGz
YlxLdn0q4u3CTC0Or05Aq3NK6eYSv68Y8CaMYEiVn92AcSCtTyfHYNMJtV8JD6ZY
7KMAEIpS/H0w9uln7y4y8uEMFzw6Dp3kM85vTPUzDQI+x2G5azR0w91lP0I0eU9Y
jWo3PwdCOe1HrR190LbbV/zNm2+ZWfQldCHCgDUhlDGJU2/ZM3KlK8vDa/rYKzQ/
mX28tJTMG0EIdwsXaPhYlrBDDwstpX/pWgCFyjq4CCCEOjjHuHU+sUYgJLawrOvF
zQOUnzOZN96+684qhp4Pf8HIKjLe0lcB4lLJOXZOCuBO2J1GVFI6lmOeC5eW2WWI
F5Ti3EvdY95yci8bKhJ5R/Hy1dY7u9wusJm7A1efMZjE3X75SZh7GLTxDl0I8l+7
JS4E6m6Axog0FZdOQvrhBB24XHWW9PdBWNr/9TW/Tbnlw3Frk5hAVFKpjv6w1ChK
fNzlbR8S8RTEn6NLQzQiYjSUZzG6QB+iTKtyoM7kAIPiWnxtDwxwFlhLkze/ZFNz
Xox+BWKUKBr0bHV3QxL2PqcFGXGU9igtnTcOh5l7IwIESMmFADxy0qYMoEiaL02M
HG851VNAWrhHOfBCQw2NmnfPN1w7r4EagdwaeuOjlE/mF+XWcbMYn9ZUvrogKHbE
VPcOdy4+DSTcgJ6aosLl8x0NR2aKf181mjflNy34ExoV6Q/IuKoAJfZqqhaotzID
755e1KtLoxm7DiBqRvrgEbEe/yhHq/QfGMqCCqxra8wXjjVCf5UigW7HvNw/JcQy
TvvtjU07/BiNOeqURtFkBYpTOFWpx7qj7fbqb46itgixpA8//dChCnNmt34BOqR5
yeeSINn9dpVrpffR3hq2MPZmTYxwwvFlMwBNS2VcFS8zsg7+ubqhen1EEuZJrh7J
XWeI89mq2WoLxMMppgf4l7v+BfE5ttalPhm/G5LFzQsafW1KknUG8Uh+6tfL0RXK
/GxpRV/oefCfUvz6MhT960x7TL2d7IP0oEDgM8oY3EDqMGgZSpwt5KxA4npEi1/I
cbaHm3PCHNyE3UAS6D3HxCIzeaxjdcG95ohjd9NmahMugwBpacciFkvneJr+IO08
KjVCq4otlmyme12RXroC6rJ/gkaAn7IsBY/GcVihVHDAJgaIy8k0AxUakCrWbv17
w+1UoLP7VWQlCb+cf6BlpklGSoNFv2ztWBR6/AMq/PYQvxy8HFRJ2jPozOyE3ckb
Y1jLbAam0bzvdfhjgR1zbIq+sV0PWOuRYHJJsXi2nn+X1repwhF4BgrzS9PJaBYD
f3ZFbHZg90qf2i4xRu0FUZ5yZFViN7fNE69e06EtryQZjQx8uJ37yYvMVo0dPnPE
+UO7Y3LfzjceqVeoMp8Lfqs5j2R7WO95W3hcr6iUnRoVLk3BjtB+Uf+bXMmBH34J
OLrYCWtPG7hhz/2kF92P70j68sIevixNojSQ3mCdpiLECu45UcJNFpLHaiu6AXAi
gOptVp34GKO/k/uX+c3UI0oR1H/jTspJdMFDVLlTlVVU8ioLDw+TPQUTTBnt0UPc
DDP3s/zRYPGL4jnM5ZozQJD3MN0gBltAsxPNuz/RNWWS7CfJU3IotUYRzwhfYZ7c
qHI8DBSGPjB7Mgad+vG7sjeLJplgSM4QF2c9CxVz1yEumbUSHn4A2cJPJrg6OHZ1
QbN2cjAcODdBbP+Cye/2wot4Bn4/K5zUELl5cm8iEpSmxgT8gATtxtPlIIyxASep
LVDX6pAM3AkD82kGOsbHs6DdJgo54a013avp6U7nnR9v42vIZwyURyBGU5N0lKTo
87/SzB7U98qp/5SppVArvPTO8YEeCR/Oyx4Wm7EmAMJPKgZloqAgCXHLZDwheDQ3
8eHg1I3ZUH/eDYcfwTsMzfOV6rxKaBNmcbl4XQgssAZfhM8mZubhfo04XDRK/dkr
3FDh4nVEZYu+4XQ8Ir+TO/Y9XcGlyzs1ycYenU3tR5JgDKc78YIzH+YJ2wUSJyh+
vd/VEi2vJwJhoKEjIsqxTaqApEunCdKkMBSoJpom2Bk+dGKyUZn5muTwVl+isnSP
scIHJp5Z9EKqIzyC1KTNGpaoI63BRWFovRZgQKn22y2gP19vL9fqoq4Rw/Upfy+B
uwd5h1Q3UVCwrp8mdsMOS/e05RdzY631aG8v7aePLPOpGZs0Vfyn5bY/eMKyWMdb
s75LHEvp27yVXyh7/FOTiKH4VIn0goA3Lv5FQiY6KLJwXVXF0zowNjJmuXeByWPi
yLxdFajZSrfZF+p6bC2lu81LB/JA6lT1iexkPe//PyrhjNUba1bzGAgoJkiwKtlF
mQlLNUAnMm7rFNMEXS9dY4yNPDlzyOe1bMcDdabktgokiOKboY/pNlYi4EIaoHZQ
wgy9/4CChpHiI6jhHZXrGSSgjpAFZBwxflUy0u5OhVN5QL4h6odi6T9wW55sDfFm
ddClAnM8rGC/fWOAFjsZK+/kcPu1puQ6UJGp1k4gBGYjwo1xi/61dzbvp+LvMSuT
YA85CuJy+CxNcnAPXuu87ffRJsikjouX0zyCe6bFK+s+pRsDYY/oBI+HGRk44OWV
G7Ejtp5cQfZ83sCHWtuHltf6MeH0R4LU/PfHkvaPS4Y24ICHEXDW8jIJWW76Hldr
kPZ3gDAklxvUtbAuV9m8fm3Xb4Njqs1LG97W46qCEmK5Eu0AS+cgH+zvXoyBfkpm
uOB436ds9zn76M59aD5dTn3XWrqdHv14l3MFwRM8GBUSiAmE75hyoHK719/SmQMo
bhg7bE76qKlTSJfeSyKYgcutqkjOWGBAdeBLS1bhRhDlM/cqLdTU3V4PlEUOF7nP
4d8FNvUV/4zdu4sQq4HJ4f5JfrXxCupeMNyB+nDfor3i9Z7V1UKcwChN1hXwN96t
O5MZgtECv10BYfSrr2Y9N6PsSFdsrPPTF/c67I3ooZfFH6QthqN5fgmog0lG/JPu
zsRRIOZs9B+wTBS3wCmskkNYk1tp85Vg6cLVhxDxEVo9jphyYs349jYcC4A9ILmd
yc3nZp/8e10El3x0V/8sx2oxB4RlkQLMPKg78WNPDDIpmz66Yu1dTLN3Kgs7bISd
Lt6B2c0MkmhoWuLAte0PB3HszTvcUrCoXSJ4MT8foCpVQFzjM3pWLQbdZLTb/eS8
C8CdVqZFV/FxTvvCMkuvnKHkBlT4WS00mxR+XcSfH0hIDsM7B0aAgbVrtpunGYlo
E98CojbeUSxy6omPrI8QepTl5cptf2JsN+XYRd2SfHLNxQhSyYqhZnNUHUK/h8gs
Zmh42EmJ13ugIfy6sCWMjsRlvjpcrybePWaVaESQkS1IbFKKdwJcYmRfdnFkaL9D
BHo+/r+V/VHZztZwRIJld68PbXawdqkdRPa89d3UfJOR6KXzMYrh/swveIBGBTfN
qgmRZ6NTrrdTwjww/Kve0FrzWr525VU3O7drtBQa6MDcbRKirPN+QY8Q6Gz8nTw0
OSgFKEJQOP2WnH9mtHxemiNW3k+FmC8rqx8r0dGp5kwFu58/9gc31cMvn0Y9RSC6
jnrbRB02srDiykVfURwGePdlz8/R/9pLZ9PYs0c2lFRKtYUvvu6WE53l9kc/rAJY
GMtArnsIcE9JDH8Dzkr1QhaxIOrKAfyHBmgYHWA6MISGp72s9cKiWdM7DNkzO4OU
/mTwrgUJ/EDEpiGIIOkZq/8FlzI9edpTsq0jGfkQuE7pLJYz/I4vgF29jgGycqBK
jKfw5scC2swO08uSOolG+A7pxkDmAa67ML8M6TtiffEbwsD2fKVBZfvbJkQFCBW6
YiHASO0KI6PrDWUWl7ghMVEmsu3q0VvQKbn098z9no1EIBCXDFgn4U0K8K8+Mrll
i5qsUy9m3b3G9cjvFrO4TSi5wHYdM8nLban1nFgVM6Q+TqwQclZsb71gbUhRcK8W
`pragma protect end_protected
