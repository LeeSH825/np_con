-- avlm_avls_1x1.vhd

-- Generated using ACDS version 21.1 842

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity avlm_avls_1x1 is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity avlm_avls_1x1;

architecture rtl of avlm_avls_1x1 is
	component altera_avalon_mm_master_bfm is
		generic (
			AV_ADDRESS_W               : integer := 32;
			AV_SYMBOL_W                : integer := 8;
			AV_NUMSYMBOLS              : integer := 4;
			AV_BURSTCOUNT_W            : integer := 3;
			AV_READRESPONSE_W          : integer := 8;
			AV_WRITERESPONSE_W         : integer := 8;
			USE_READ                   : integer := 1;
			USE_WRITE                  : integer := 1;
			USE_ADDRESS                : integer := 1;
			USE_BYTE_ENABLE            : integer := 1;
			USE_BURSTCOUNT             : integer := 1;
			USE_READ_DATA              : integer := 1;
			USE_READ_DATA_VALID        : integer := 1;
			USE_WRITE_DATA             : integer := 1;
			USE_BEGIN_TRANSFER         : integer := 0;
			USE_BEGIN_BURST_TRANSFER   : integer := 0;
			USE_WAIT_REQUEST           : integer := 1;
			USE_TRANSACTIONID          : integer := 0;
			USE_WRITERESPONSE          : integer := 0;
			USE_READRESPONSE           : integer := 0;
			USE_CLKEN                  : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR : integer := 1;
			AV_BURST_LINEWRAP          : integer := 1;
			AV_BURST_BNDR_ONLY         : integer := 1;
			AV_MAX_PENDING_READS       : integer := 0;
			AV_MAX_PENDING_WRITES      : integer := 0;
			AV_FIX_READ_LATENCY        : integer := 1;
			AV_READ_WAIT_TIME          : integer := 1;
			AV_WRITE_WAIT_TIME         : integer := 0;
			REGISTER_WAITREQUEST       : integer := 0;
			AV_REGISTERINCOMINGSIGNALS : integer := 0;
			VHDL_ID                    : integer := 0
		);
		port (
			clk                    : in  std_logic                     := 'X';             -- clk
			reset                  : in  std_logic                     := 'X';             -- reset
			avm_address            : out std_logic_vector(31 downto 0);                    -- address
			avm_burstcount         : out std_logic_vector(3 downto 0);                     -- burstcount
			avm_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			avm_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			avm_write              : out std_logic;                                        -- write
			avm_read               : out std_logic;                                        -- read
			avm_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			avm_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			avm_begintransfer      : out std_logic;                                        -- begintransfer
			avm_beginbursttransfer : out std_logic;                                        -- beginbursttransfer
			avm_arbiterlock        : out std_logic;                                        -- arbiterlock
			avm_lock               : out std_logic;                                        -- lock
			avm_debugaccess        : out std_logic;                                        -- debugaccess
			avm_transactionid      : out std_logic_vector(7 downto 0);                     -- transactionid
			avm_readid             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readid
			avm_writeid            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writeid
			avm_clken              : out std_logic;                                        -- clken
			avm_response           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			avm_writeresponsevalid : in  std_logic                     := 'X';             -- writeresponsevalid
			avm_readresponse       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readresponse
			avm_writeresponse      : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- writeresponse
		);
	end component altera_avalon_mm_master_bfm;

	component addr_slave is
		generic (
			ADDRESS_WIDTH : integer := 12;
			BURST_WIDTH   : integer := 4;
			BYTE_WIDTH    : integer := 4;
			DATA_WIDTH    : integer := 32
		);
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			avs_s0_address     : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			avs_s0_waitrequest : out std_logic;                                        -- waitrequest
			avs_s0_burstcount  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			avs_s0_byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_s0_write       : in  std_logic                     := 'X';             -- write
			avs_s0_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avm_m0_address     : out std_logic_vector(11 downto 0);                    -- address
			avm_m0_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			avm_m0_burstcount  : out std_logic_vector(3 downto 0);                     -- burstcount
			avm_m0_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			avm_m0_write       : out std_logic;                                        -- write
			avm_m0_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			rst                : in  std_logic                     := 'X'              -- reset
		);
	end component addr_slave;

	component altera_avalon_mm_slave_bfm is
		generic (
			AV_ADDRESS_W               : integer := 32;
			AV_SYMBOL_W                : integer := 8;
			AV_NUMSYMBOLS              : integer := 4;
			AV_BURSTCOUNT_W            : integer := 3;
			AV_READRESPONSE_W          : integer := 8;
			AV_WRITERESPONSE_W         : integer := 8;
			USE_READ                   : integer := 1;
			USE_WRITE                  : integer := 1;
			USE_ADDRESS                : integer := 1;
			USE_BYTE_ENABLE            : integer := 1;
			USE_BURSTCOUNT             : integer := 1;
			USE_READ_DATA              : integer := 1;
			USE_READ_DATA_VALID        : integer := 1;
			USE_WRITE_DATA             : integer := 1;
			USE_BEGIN_TRANSFER         : integer := 0;
			USE_BEGIN_BURST_TRANSFER   : integer := 0;
			USE_WAIT_REQUEST           : integer := 1;
			USE_TRANSACTIONID          : integer := 0;
			USE_WRITERESPONSE          : integer := 0;
			USE_READRESPONSE           : integer := 0;
			USE_CLKEN                  : integer := 0;
			AV_BURST_LINEWRAP          : integer := 1;
			AV_BURST_BNDR_ONLY         : integer := 1;
			AV_MAX_PENDING_READS       : integer := 1;
			AV_MAX_PENDING_WRITES      : integer := 0;
			AV_FIX_READ_LATENCY        : integer := 0;
			AV_READ_WAIT_TIME          : integer := 1;
			AV_WRITE_WAIT_TIME         : integer := 0;
			REGISTER_WAITREQUEST       : integer := 0;
			AV_REGISTERINCOMINGSIGNALS : integer := 0;
			VHDL_ID                    : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			avs_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_burstcount           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			avs_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			avs_address              : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			avs_waitrequest          : out std_logic;                                        -- waitrequest
			avs_write                : in  std_logic                     := 'X';             -- write
			avs_read                 : in  std_logic                     := 'X';             -- read
			avs_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_readdatavalid        : out std_logic;                                        -- readdatavalid
			avs_begintransfer        : in  std_logic                     := 'X';             -- begintransfer
			avs_beginbursttransfer   : in  std_logic                     := 'X';             -- beginbursttransfer
			avs_arbiterlock          : in  std_logic                     := 'X';             -- arbiterlock
			avs_lock                 : in  std_logic                     := 'X';             -- lock
			avs_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			avs_transactionid        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- transactionid
			avs_readid               : out std_logic_vector(7 downto 0);                     -- readid
			avs_writeid              : out std_logic_vector(7 downto 0);                     -- writeid
			avs_clken                : in  std_logic                     := 'X';             -- clken
			avs_response             : out std_logic_vector(1 downto 0);                     -- response
			avs_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			avs_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			avs_readresponse         : out std_logic_vector(7 downto 0);                     -- readresponse
			avs_writeresponse        : out std_logic_vector(7 downto 0)                      -- writeresponse
		);
	end component altera_avalon_mm_slave_bfm;

	component avlm_avls_1x1_mm_interconnect_0 is
		port (
			clk_clk_clk                                    : in  std_logic                     := 'X';             -- clk
			master_0_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			master_0_m0_address                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			master_0_m0_waitrequest                        : out std_logic;                                        -- waitrequest
			master_0_m0_burstcount                         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			master_0_m0_byteenable                         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			master_0_m0_read                               : in  std_logic                     := 'X';             -- read
			master_0_m0_readdata                           : out std_logic_vector(31 downto 0);                    -- readdata
			master_0_m0_readdatavalid                      : out std_logic;                                        -- readdatavalid
			master_0_m0_write                              : in  std_logic                     := 'X';             -- write
			master_0_m0_writedata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			monitor_0_s0_address                           : out std_logic_vector(11 downto 0);                    -- address
			monitor_0_s0_write                             : out std_logic;                                        -- write
			monitor_0_s0_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			monitor_0_s0_burstcount                        : out std_logic_vector(3 downto 0);                     -- burstcount
			monitor_0_s0_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			monitor_0_s0_waitrequest                       : in  std_logic                     := 'X'              -- waitrequest
		);
	end component avlm_avls_1x1_mm_interconnect_0;

	component avlm_avls_1x1_mm_interconnect_1 is
		port (
			clk_clk_clk                                      : in  std_logic                     := 'X';             -- clk
			monitor_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			monitor_0_m0_address                             : in  std_logic_vector(11 downto 0) := (others => 'X'); -- address
			monitor_0_m0_waitrequest                         : out std_logic;                                        -- waitrequest
			monitor_0_m0_burstcount                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			monitor_0_m0_byteenable                          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			monitor_0_m0_write                               : in  std_logic                     := 'X';             -- write
			monitor_0_m0_writedata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_0_s0_address                               : out std_logic_vector(11 downto 0);                    -- address
			slave_0_s0_write                                 : out std_logic;                                        -- write
			slave_0_s0_read                                  : out std_logic;                                        -- read
			slave_0_s0_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			slave_0_s0_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			slave_0_s0_burstcount                            : out std_logic_vector(3 downto 0);                     -- burstcount
			slave_0_s0_byteenable                            : out std_logic_vector(3 downto 0);                     -- byteenable
			slave_0_s0_readdatavalid                         : in  std_logic                     := 'X';             -- readdatavalid
			slave_0_s0_waitrequest                           : in  std_logic                     := 'X'              -- waitrequest
		);
	end component avlm_avls_1x1_mm_interconnect_1;

	signal master_0_m0_readdata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:master_0_m0_readdata -> master_0:avm_readdata
	signal master_0_m0_waitrequest                    : std_logic;                     -- mm_interconnect_0:master_0_m0_waitrequest -> master_0:avm_waitrequest
	signal master_0_m0_address                        : std_logic_vector(31 downto 0); -- master_0:avm_address -> mm_interconnect_0:master_0_m0_address
	signal master_0_m0_read                           : std_logic;                     -- master_0:avm_read -> mm_interconnect_0:master_0_m0_read
	signal master_0_m0_byteenable                     : std_logic_vector(3 downto 0);  -- master_0:avm_byteenable -> mm_interconnect_0:master_0_m0_byteenable
	signal master_0_m0_readdatavalid                  : std_logic;                     -- mm_interconnect_0:master_0_m0_readdatavalid -> master_0:avm_readdatavalid
	signal master_0_m0_writedata                      : std_logic_vector(31 downto 0); -- master_0:avm_writedata -> mm_interconnect_0:master_0_m0_writedata
	signal master_0_m0_write                          : std_logic;                     -- master_0:avm_write -> mm_interconnect_0:master_0_m0_write
	signal master_0_m0_burstcount                     : std_logic_vector(3 downto 0);  -- master_0:avm_burstcount -> mm_interconnect_0:master_0_m0_burstcount
	signal mm_interconnect_0_monitor_0_s0_waitrequest : std_logic;                     -- monitor_0:avs_s0_waitrequest -> mm_interconnect_0:monitor_0_s0_waitrequest
	signal mm_interconnect_0_monitor_0_s0_address     : std_logic_vector(11 downto 0); -- mm_interconnect_0:monitor_0_s0_address -> monitor_0:avs_s0_address
	signal mm_interconnect_0_monitor_0_s0_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:monitor_0_s0_byteenable -> monitor_0:avs_s0_byteenable
	signal mm_interconnect_0_monitor_0_s0_write       : std_logic;                     -- mm_interconnect_0:monitor_0_s0_write -> monitor_0:avs_s0_write
	signal mm_interconnect_0_monitor_0_s0_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:monitor_0_s0_writedata -> monitor_0:avs_s0_writedata
	signal mm_interconnect_0_monitor_0_s0_burstcount  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:monitor_0_s0_burstcount -> monitor_0:avs_s0_burstcount
	signal monitor_0_m0_waitrequest                   : std_logic;                     -- mm_interconnect_1:monitor_0_m0_waitrequest -> monitor_0:avm_m0_waitrequest
	signal monitor_0_m0_address                       : std_logic_vector(11 downto 0); -- monitor_0:avm_m0_address -> mm_interconnect_1:monitor_0_m0_address
	signal monitor_0_m0_byteenable                    : std_logic_vector(3 downto 0);  -- monitor_0:avm_m0_byteenable -> mm_interconnect_1:monitor_0_m0_byteenable
	signal monitor_0_m0_write                         : std_logic;                     -- monitor_0:avm_m0_write -> mm_interconnect_1:monitor_0_m0_write
	signal monitor_0_m0_writedata                     : std_logic_vector(31 downto 0); -- monitor_0:avm_m0_writedata -> mm_interconnect_1:monitor_0_m0_writedata
	signal monitor_0_m0_burstcount                    : std_logic_vector(3 downto 0);  -- monitor_0:avm_m0_burstcount -> mm_interconnect_1:monitor_0_m0_burstcount
	signal mm_interconnect_1_slave_0_s0_readdata      : std_logic_vector(31 downto 0); -- slave_0:avs_readdata -> mm_interconnect_1:slave_0_s0_readdata
	signal mm_interconnect_1_slave_0_s0_waitrequest   : std_logic;                     -- slave_0:avs_waitrequest -> mm_interconnect_1:slave_0_s0_waitrequest
	signal mm_interconnect_1_slave_0_s0_address       : std_logic_vector(11 downto 0); -- mm_interconnect_1:slave_0_s0_address -> slave_0:avs_address
	signal mm_interconnect_1_slave_0_s0_read          : std_logic;                     -- mm_interconnect_1:slave_0_s0_read -> slave_0:avs_read
	signal mm_interconnect_1_slave_0_s0_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_1:slave_0_s0_byteenable -> slave_0:avs_byteenable
	signal mm_interconnect_1_slave_0_s0_readdatavalid : std_logic;                     -- slave_0:avs_readdatavalid -> mm_interconnect_1:slave_0_s0_readdatavalid
	signal mm_interconnect_1_slave_0_s0_write         : std_logic;                     -- mm_interconnect_1:slave_0_s0_write -> slave_0:avs_write
	signal mm_interconnect_1_slave_0_s0_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_1:slave_0_s0_writedata -> slave_0:avs_writedata
	signal mm_interconnect_1_slave_0_s0_burstcount    : std_logic_vector(3 downto 0);  -- mm_interconnect_1:slave_0_s0_burstcount -> slave_0:avs_burstcount
	signal reset_reset_n_ports_inv                    : std_logic;                     -- reset_reset_n:inv -> [master_0:reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:monitor_0_reset_sink_reset_bridge_in_reset_reset, monitor_0:rst, slave_0:reset]

begin

	master_0 : component altera_avalon_mm_master_bfm
		generic map (
			AV_ADDRESS_W               => 32,
			AV_SYMBOL_W                => 8,
			AV_NUMSYMBOLS              => 4,
			AV_BURSTCOUNT_W            => 4,
			AV_READRESPONSE_W          => 8,
			AV_WRITERESPONSE_W         => 8,
			USE_READ                   => 1,
			USE_WRITE                  => 1,
			USE_ADDRESS                => 1,
			USE_BYTE_ENABLE            => 1,
			USE_BURSTCOUNT             => 1,
			USE_READ_DATA              => 1,
			USE_READ_DATA_VALID        => 1,
			USE_WRITE_DATA             => 1,
			USE_BEGIN_TRANSFER         => 0,
			USE_BEGIN_BURST_TRANSFER   => 0,
			USE_WAIT_REQUEST           => 1,
			USE_TRANSACTIONID          => 0,
			USE_WRITERESPONSE          => 0,
			USE_READRESPONSE           => 0,
			USE_CLKEN                  => 0,
			AV_CONSTANT_BURST_BEHAVIOR => 1,
			AV_BURST_LINEWRAP          => 0,
			AV_BURST_BNDR_ONLY         => 0,
			AV_MAX_PENDING_READS       => 8,
			AV_MAX_PENDING_WRITES      => 0,
			AV_FIX_READ_LATENCY        => 0,
			AV_READ_WAIT_TIME          => 1,
			AV_WRITE_WAIT_TIME         => 0,
			REGISTER_WAITREQUEST       => 0,
			AV_REGISTERINCOMINGSIGNALS => 0,
			VHDL_ID                    => 0
		)
		port map (
			clk                    => clk_clk,                   --       clk.clk
			reset                  => reset_reset_n_ports_inv,   -- clk_reset.reset
			avm_address            => master_0_m0_address,       --        m0.address
			avm_burstcount         => master_0_m0_burstcount,    --          .burstcount
			avm_readdata           => master_0_m0_readdata,      --          .readdata
			avm_writedata          => master_0_m0_writedata,     --          .writedata
			avm_waitrequest        => master_0_m0_waitrequest,   --          .waitrequest
			avm_write              => master_0_m0_write,         --          .write
			avm_read               => master_0_m0_read,          --          .read
			avm_byteenable         => master_0_m0_byteenable,    --          .byteenable
			avm_readdatavalid      => master_0_m0_readdatavalid, --          .readdatavalid
			avm_begintransfer      => open,                      -- (terminated)
			avm_beginbursttransfer => open,                      -- (terminated)
			avm_arbiterlock        => open,                      -- (terminated)
			avm_lock               => open,                      -- (terminated)
			avm_debugaccess        => open,                      -- (terminated)
			avm_transactionid      => open,                      -- (terminated)
			avm_readid             => "00000000",                -- (terminated)
			avm_writeid            => "00000000",                -- (terminated)
			avm_clken              => open,                      -- (terminated)
			avm_response           => "00",                      -- (terminated)
			avm_writeresponsevalid => '0',                       -- (terminated)
			avm_readresponse       => "00000000",                -- (terminated)
			avm_writeresponse      => "00000000"                 -- (terminated)
		);

	monitor_0 : component addr_slave
		generic map (
			ADDRESS_WIDTH => 12,
			BURST_WIDTH   => 4,
			BYTE_WIDTH    => 4,
			DATA_WIDTH    => 32
		)
		port map (
			clk                => clk_clk,                                    --      clock.clk
			avs_s0_address     => mm_interconnect_0_monitor_0_s0_address,     --         s0.address
			avs_s0_waitrequest => mm_interconnect_0_monitor_0_s0_waitrequest, --           .waitrequest
			avs_s0_burstcount  => mm_interconnect_0_monitor_0_s0_burstcount,  --           .burstcount
			avs_s0_byteenable  => mm_interconnect_0_monitor_0_s0_byteenable,  --           .byteenable
			avs_s0_write       => mm_interconnect_0_monitor_0_s0_write,       --           .write
			avs_s0_writedata   => mm_interconnect_0_monitor_0_s0_writedata,   --           .writedata
			avm_m0_address     => monitor_0_m0_address,                       --         m0.address
			avm_m0_waitrequest => monitor_0_m0_waitrequest,                   --           .waitrequest
			avm_m0_burstcount  => monitor_0_m0_burstcount,                    --           .burstcount
			avm_m0_byteenable  => monitor_0_m0_byteenable,                    --           .byteenable
			avm_m0_write       => monitor_0_m0_write,                         --           .write
			avm_m0_writedata   => monitor_0_m0_writedata,                     --           .writedata
			rst                => reset_reset_n_ports_inv                     -- reset_sink.reset
		);

	slave_0 : component altera_avalon_mm_slave_bfm
		generic map (
			AV_ADDRESS_W               => 12,
			AV_SYMBOL_W                => 8,
			AV_NUMSYMBOLS              => 4,
			AV_BURSTCOUNT_W            => 4,
			AV_READRESPONSE_W          => 8,
			AV_WRITERESPONSE_W         => 8,
			USE_READ                   => 1,
			USE_WRITE                  => 1,
			USE_ADDRESS                => 1,
			USE_BYTE_ENABLE            => 1,
			USE_BURSTCOUNT             => 1,
			USE_READ_DATA              => 1,
			USE_READ_DATA_VALID        => 1,
			USE_WRITE_DATA             => 1,
			USE_BEGIN_TRANSFER         => 0,
			USE_BEGIN_BURST_TRANSFER   => 0,
			USE_WAIT_REQUEST           => 1,
			USE_TRANSACTIONID          => 0,
			USE_WRITERESPONSE          => 0,
			USE_READRESPONSE           => 0,
			USE_CLKEN                  => 0,
			AV_BURST_LINEWRAP          => 0,
			AV_BURST_BNDR_ONLY         => 0,
			AV_MAX_PENDING_READS       => 1,
			AV_MAX_PENDING_WRITES      => 0,
			AV_FIX_READ_LATENCY        => 0,
			AV_READ_WAIT_TIME          => 1,
			AV_WRITE_WAIT_TIME         => 0,
			REGISTER_WAITREQUEST       => 0,
			AV_REGISTERINCOMINGSIGNALS => 0,
			VHDL_ID                    => 0
		)
		port map (
			clk                      => clk_clk,                                    --       clk.clk
			reset                    => reset_reset_n_ports_inv,                    -- clk_reset.reset
			avs_writedata            => mm_interconnect_1_slave_0_s0_writedata,     --        s0.writedata
			avs_burstcount           => mm_interconnect_1_slave_0_s0_burstcount,    --          .burstcount
			avs_readdata             => mm_interconnect_1_slave_0_s0_readdata,      --          .readdata
			avs_address              => mm_interconnect_1_slave_0_s0_address,       --          .address
			avs_waitrequest          => mm_interconnect_1_slave_0_s0_waitrequest,   --          .waitrequest
			avs_write                => mm_interconnect_1_slave_0_s0_write,         --          .write
			avs_read                 => mm_interconnect_1_slave_0_s0_read,          --          .read
			avs_byteenable           => mm_interconnect_1_slave_0_s0_byteenable,    --          .byteenable
			avs_readdatavalid        => mm_interconnect_1_slave_0_s0_readdatavalid, --          .readdatavalid
			avs_begintransfer        => '0',                                        -- (terminated)
			avs_beginbursttransfer   => '0',                                        -- (terminated)
			avs_arbiterlock          => '0',                                        -- (terminated)
			avs_lock                 => '0',                                        -- (terminated)
			avs_debugaccess          => '0',                                        -- (terminated)
			avs_transactionid        => "00000000",                                 -- (terminated)
			avs_readid               => open,                                       -- (terminated)
			avs_writeid              => open,                                       -- (terminated)
			avs_clken                => '1',                                        -- (terminated)
			avs_response             => open,                                       -- (terminated)
			avs_writeresponserequest => '0',                                        -- (terminated)
			avs_writeresponsevalid   => open,                                       -- (terminated)
			avs_readresponse         => open,                                       -- (terminated)
			avs_writeresponse        => open                                        -- (terminated)
		);

	mm_interconnect_0 : component avlm_avls_1x1_mm_interconnect_0
		port map (
			clk_clk_clk                                    => clk_clk,                                    --                                  clk_clk.clk
			master_0_clk_reset_reset_bridge_in_reset_reset => reset_reset_n_ports_inv,                    -- master_0_clk_reset_reset_bridge_in_reset.reset
			master_0_m0_address                            => master_0_m0_address,                        --                              master_0_m0.address
			master_0_m0_waitrequest                        => master_0_m0_waitrequest,                    --                                         .waitrequest
			master_0_m0_burstcount                         => master_0_m0_burstcount,                     --                                         .burstcount
			master_0_m0_byteenable                         => master_0_m0_byteenable,                     --                                         .byteenable
			master_0_m0_read                               => master_0_m0_read,                           --                                         .read
			master_0_m0_readdata                           => master_0_m0_readdata,                       --                                         .readdata
			master_0_m0_readdatavalid                      => master_0_m0_readdatavalid,                  --                                         .readdatavalid
			master_0_m0_write                              => master_0_m0_write,                          --                                         .write
			master_0_m0_writedata                          => master_0_m0_writedata,                      --                                         .writedata
			monitor_0_s0_address                           => mm_interconnect_0_monitor_0_s0_address,     --                             monitor_0_s0.address
			monitor_0_s0_write                             => mm_interconnect_0_monitor_0_s0_write,       --                                         .write
			monitor_0_s0_writedata                         => mm_interconnect_0_monitor_0_s0_writedata,   --                                         .writedata
			monitor_0_s0_burstcount                        => mm_interconnect_0_monitor_0_s0_burstcount,  --                                         .burstcount
			monitor_0_s0_byteenable                        => mm_interconnect_0_monitor_0_s0_byteenable,  --                                         .byteenable
			monitor_0_s0_waitrequest                       => mm_interconnect_0_monitor_0_s0_waitrequest  --                                         .waitrequest
		);

	mm_interconnect_1 : component avlm_avls_1x1_mm_interconnect_1
		port map (
			clk_clk_clk                                      => clk_clk,                                    --                                    clk_clk.clk
			monitor_0_reset_sink_reset_bridge_in_reset_reset => reset_reset_n_ports_inv,                    -- monitor_0_reset_sink_reset_bridge_in_reset.reset
			monitor_0_m0_address                             => monitor_0_m0_address,                       --                               monitor_0_m0.address
			monitor_0_m0_waitrequest                         => monitor_0_m0_waitrequest,                   --                                           .waitrequest
			monitor_0_m0_burstcount                          => monitor_0_m0_burstcount,                    --                                           .burstcount
			monitor_0_m0_byteenable                          => monitor_0_m0_byteenable,                    --                                           .byteenable
			monitor_0_m0_write                               => monitor_0_m0_write,                         --                                           .write
			monitor_0_m0_writedata                           => monitor_0_m0_writedata,                     --                                           .writedata
			slave_0_s0_address                               => mm_interconnect_1_slave_0_s0_address,       --                                 slave_0_s0.address
			slave_0_s0_write                                 => mm_interconnect_1_slave_0_s0_write,         --                                           .write
			slave_0_s0_read                                  => mm_interconnect_1_slave_0_s0_read,          --                                           .read
			slave_0_s0_readdata                              => mm_interconnect_1_slave_0_s0_readdata,      --                                           .readdata
			slave_0_s0_writedata                             => mm_interconnect_1_slave_0_s0_writedata,     --                                           .writedata
			slave_0_s0_burstcount                            => mm_interconnect_1_slave_0_s0_burstcount,    --                                           .burstcount
			slave_0_s0_byteenable                            => mm_interconnect_1_slave_0_s0_byteenable,    --                                           .byteenable
			slave_0_s0_readdatavalid                         => mm_interconnect_1_slave_0_s0_readdatavalid, --                                           .readdatavalid
			slave_0_s0_waitrequest                           => mm_interconnect_1_slave_0_s0_waitrequest    --                                           .waitrequest
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

end architecture rtl; -- of avlm_avls_1x1
