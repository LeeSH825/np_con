library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package PROPERTIES_PACK is
	
	constant DATA_WIDTH		: integer			:= 8;
	constant ADDR_WIDTH		: integer			:= 2;

end package PROPERTIES_PACK;

-- package body PROPERTIES_PACK is
-- 	generic map (DATA_WIDTH => 8,
-- 				ADDR_WIDTH => 2)
	
	
-- end package body PROPERTIES_PACK;