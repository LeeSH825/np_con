`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZqR8iE2VxBNRC2MT9xxRGq7yTJu/d5+TOkxBWtQriw2UfbW/+7M8kpXXhSVuNZ+2
JapbdFvg78vWXDDI+DPMT4WLGe/9f4PmZ+ws/zPC3VNqNU/zFqfwS+5HCj00JoGP
otgFXBIUf2v5fd6gOTk7OErfDduafWzV5DCR+yOobho=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57024)
9uoczLBD+bcaRIZ70b2J3mIoAuH6RjD/Jn2veIOyDIbAL4fGA563H93zmv2VGlHB
mAuFlj+wFng9IfXttDRa9hhrx826IvhpmSgSzdatnvrHR/XED9zRxxVBdlC+F1wu
5bdj1WNLySBsRoPm7l4os6lyiUYFV6JGVe2RpbxLKGDQZeH/il4QqfmCL0toEp1e
PflSuX56Nl1AUSmx5f7DrEUonTrcOo31H6GNNCz2OFFgyatGcVOoGRYCfJwrg/xJ
QdeAeeszP+02yv6Civ5DdxeNv1jUo8jkVCy2MxbItfIRgyMiVnTrcxmD6V5TIMzD
cvCaT3ncGAol4Yk447GUOJOuge28pj+PbcE+ZBlWZXzqbFkYT5BcNq7TNqwUsnGa
754o2LrIAvoz3PItGh29dy8/Sm6V2qQxZJrokNdN0WqHQWzIiVY/LjZquc7Cjx21
pkK9wiNXlQEKT2W4WVVGffWfL5WNVD/6IIPl8ViBU37dBp8WojKubTfOy69ROy2z
2ar7qDwd7x9gp3QwcZXdkKY+TZvxPkEAOK2EW6bdAkFrQK3WlXMHiil4yHfhQhwL
WhNuUOrSfI4VHihSodr2AZGFTlZk7fdk7fn7nKIRe+FkHvRlS5Xu1BF84GGc/HBs
0++4y31KqO/Cwa2vBWVSaIylmK+zWLKULN8X7+7p5wWDji8dLtMKcpj7639lAADt
CUWHj/ZjMaoyJE21fVoU++NLZAR4IIJNzuqvtJ5WEnkGp6FIjaNZmaozQl9Xc5un
zUeUTHo6ofGvD8ZK32DfPxhXLzy5qMThDo3Ovxyx7wcZTEKEcUpNY+vPBIrwrGzI
fuM+NshUXMqeq2ppn9w7romvNMVpcX0M1CHvQHrxrfHnyiSVQa+V+q/jTrABMBvf
H/KV486LuUZ8XWvgyhwLHWACGkvZuX/A7adSADbcWpv5B9A4tL2Lyb6g09aytkND
ZoNj14kMRo1SP13NpbORI7+bF/k+BMfJ9YfY/NQyeyfz1GBFcOYDC85bPN8/QQ6U
Pq7EBdgDuAzipYSBRvU1UZXJsi6AcQLg2SBH+IW3Av9jVgiWtSeCxFIWS7KZYUml
XxfWjxavJTTf64QJfA6gXa07gMG0T6bvANwOT1453hWVyYcAJn3YQcldt105kvJP
pEuKOHe3FPEnMfqk3OlTalSB5qQT3zxPGK2d4QV060Ph+BfVULF/vSubHGEV2MLT
AqgRTgfiV6jHM0HcbGgeznlky9ciVaaChAK1RS/qEZAA0ga8eeoUDdOG34ei9FFB
KuSgRy9n7lUAlWYH3xWgF67yLmRgcMwNLr62BXZp70EOjsqOtr4fjuY/BdXZGgBF
TOWlvgsoXk5OCAa9mgxVnXtwW0+SYUqgcWUamQ9C8d3/x1rP3Mmsi8/AgSxpPIWr
0bp1jX2b+2ExmDzGdtR86+fFuaE07o8qT+cVEDZo+700aajaRNchFs68iSrzXN+U
42kOEZhEqa3LgVWkDr0Jnmm+K+z0gUqOA6Qr5BbJ/LLK6vDdvWT+xa7fvVZ0iZuV
Z0w3Sura+t/XX0pPy48Ly7O70RIKfiY64qDOAz6AVaK6w/LaW+dVRqCLjgMeinm8
nj9N/c8yhIfque2FIjshI+muIMDStBrXAQvzA946UrQvq6b28XAQrfBnTPed0r8b
nC/vwk+62QUDlwaxROzH9YH8LbEIptQvrd6x2eUAuX/vyvr4ax7c+/bk8AQS+RzC
f7la0dkL0I+mDe4pb0e91LlEYjJclG70r32uPn4qC/ftdCan4QeYBsteTJmde/90
XyJLOb/CFfML9XZV0ET8CJNBkmdLennFFCQbnLJ3VDrm1W0T4eixF9LtB+JadCZe
pc2YbyAgkvP8709qLtkty7eOAoCbupiNN0FiH/SL6RAUxpQo4dyovoY//DgwiPxy
MxAIVhuKucr1wt6aFM31t/NeOlG2yvruSwrKrrsqnstiiLzyUnZmB2f54k2dYKLC
et2RBIL2yCMLMdNf1H7JRA2MJVgW/17Npu0dG3L+A8iVH0JJkotXAzNIC2/UXzbv
XxTBM/X4c8DgQWLWends7x9+hMI4MsuGzghanfYd4086fOxbo55an1EskP8pLdBP
1XRCqkC3zTCcborGJDTGbvePyI8+eOVykO0Pf2pWCc4UlPB4/44qSn5q95Kzx0lB
VQBaIf0ib0NferT/wbhdpiodKPe7UPA+4qXH+7aMw3fBYpDDojgv+TZ3Lo+BD0Wp
Lix9FyMuLAtRXnWAakfe3756SS7dX4gy1OlopNRgpnHDcaXoQzoRPfovdewq1I9V
jq5z4o1vAfkIUHjQCDz+P8mEDD2tViHxFbblZGnGtIGPvfsfn9s3UHQMAT7ZLAAF
wDVGm461juEKapXenpMKHmyduEtCf40N95She4V+ctiHIBxjMRR8hifFBFx7GCwe
fNOEb9diyosPTJiaxg+LWdbD3hFcwX+BdtBfkf6IYYRnS4byD5ngFtykMC8uq+lq
17hpWxtie2uFdD62M5f8YzDehQ3Iu3HurvlgYPxuCaO1rmM007kFHP8ICaPWqQoz
fQNaJQwGd00hTzdBn2FiLfnHc9yN1SNMBQuKUDF+fG91U0fFUdWxYQWDyhYPhMB8
C/kwYJcOyKGcVMQ174ER3sZ8DH9SxCjYwdFkXe/IQWvk1tKyyNWBL2tEtYOPPUAl
2U69qZfM60hue3A5u41IxYeNQTzUFnax42haY5Y74sIObYvNvush+BrtsbzCDkW9
CY4fv2Cl4EkHCgMYE/szJPjK7r1saVWzlfdwUFAFXGxzHiKUS4NzaY0yt8TvxqGJ
hSkSls5GDAsDIXTLfdxymKp8FJgbZZIKVS3SOK104g+AwYHcseiOIGtNtRZ32Apz
CLVWMbpe0K/COV/xKncR3pJpPARYIyKDQewmoai0B+zzrz6HIPJlD5XutfJveFLI
/m6kWtkDtcv1DJGIhnRjb055iWEFqy05M4nPXxrQSv/Jxe2uSeeetN58RSTUs0le
O+krilmMFN7haIdlx4XEDDd2cVIJKQ1fYu8Lu0lgc6xgfUqPBMRjTho9x8EeTntv
IQYhbetsj+mZz3PVV+Hsusq982Ut1Q6uzaFaN+WYmrPPsoHfTnoA0tGy4UFj5WRP
7H0/aijxloOYfP15WU2Fc3RUmEzNlfJrmeAWM9uNR4lE1dwAvELvWp5gg9QnMVOU
EyrCzFzjcsv26/qMxkQuYzerxbIqQkqpAFRR902zYn7TV7mETGBlnc+s0fKFXsjf
aSC/bCits/rZTphRPZkqCWb9wXjct9vyt/9haH5JuJHH0CgcljSdjBcCD3PvSttj
K0PG7UwUXfLeg+GwvsfVIKLBuauCQeq2gYwM+PW2bhzK7rk6d+DuYeHj2hWmnNS3
+qcNHLDymk5d9iqXE4xpkMgS4dvAD9pX4DNElIExtncb8cIG/5gJPGPo1Ro/RlkT
MkzBsrCXCZdL7z5kLKlnW9eLj23IA10FXX3/jy0scVsfM0Gm96HpH/YuD/Yy1rhO
C3rZ9PJgLpS1Zbhnt9A/VYrFRSIZOmHBmFcapUXcfnnXKCos8of0lH+AkfXGxjKS
M6YVQuKlECGOLhYSLxJuJqmZLGFjz/HwAlFQ2GYSaXu/k6SE4NS1Lk+xneSIPuKF
OKFasM7UJStwZT84i/rmhG87q1xqhMBEQRcg+xHl5onB/Irpnx4tdN5gdcfZMtH3
Lsck4Sj3ySBw7qv5/tSQqrfKOs+K/PSDZnAEBHVWG7XtSpnq+lTW5UvPtWTbyRql
4C/M7qohOygaBFEUGZ0BwXPPRpJF5mEZhYlFGo6hdfWXF3c18dFJJrZeaq3xyB6G
7hTGPAuhYNPfV0wD5IbahqHggtpgIDkqnmUAMGlGztUn728QUEgGHgj5uOAmqZmp
3uzYDwdPUC3lQf/9kxTcgNG2nnay0HZU4h4U6Wgf0JZICcahroYMwET2ShKtGWb8
SLnT3Gz5YKyLSoXA0qQ9fy3E/4J9wWqB7aNxgGqir443HwHdy3UjX3JWEm6jb20y
Ql9WIXUnDNVc8T2jyDiweTxp9ZvibEgq0S4QB0gmUV6VQNyNQf8Y7yITik5x+ddm
Hap/WezuEHhB0r+59oHLpf6mvZ/tPV5dVftzXcXX8Ow+iZ1Raf2vA2UGjjg+p7mv
toOeUGT4CsCVWo8ZFeTq0SywHhTwJqdDRdaeMSKxCKr0113qAt2aA793JuM4FbZF
KZVbbgKIfqPz3t20B1EdS3n58XTrtweNvAemd6oNMmA7ktRdSGNY1qI/sJI5gY9M
RG5Cs9k9qWH6Q8zc3+4LmXFHFRbPHoFPK5PSUTIE4kzKJYEcvHwdyWhJROtLv/ib
3V6AudrVoQ0Y7a1VZb/kBtQrwKAtzlZICcWgOa2n/5E5JQ1GLwbYO/XRngH8TzXN
JLbArfxSGHBAmIT9Skrp8uA4Y6J8kDpEIgRPraJcT8r7JknTazsi9CLoQEd8RvXR
4jsmy/Mz0x5kYQZSdFYeDCOotM2nYUMFGtkFpL2cYxCMRJfdl855ASSfoEWapi6k
TUnKBShDOupaxUYVDbePjyOQxPhu6z3i6UAUcDNQWUGRiE4nBOuaXQJFBkxq9iY2
u+ew78vFHO97JWEAfyu0AfW1ONPxL8QC7kzSXNCTntvpq3C1Hylp0KjqYQiPfwMK
dae+NppxcSnD5Jt/RBCl4K2Z7DfeyQqvhWWC38H2cRVzcfF+h4ivvC8khXGE8Ljh
EWZzhk0RfE7LGJOfw23eBEJOvaZkZHlI4sO+0go28S8lOT/+EQmpbt4CBKZPeuWR
n+mvsxJqPBIXJQSiN7SHzbXaMilOIU4mK1wuFi2Td22ne5hFwXh9QEI8OSOlBTeo
kh2GK+jojMzS6df1gZAMpIXBkX/kuKZCtzSLCJsrun4zXb4pa0kk2YHsE8Q1juqm
Lcwl6JUrferhGXKwrANuTFSC4FO/GqiJWNv7cpqQVxkS2ojWzvTz3OV9LJXh32j2
AF4KxVXVxgmPn84LGHa64HmJfTC30UprQ8oK8BHNNhl7fx0dUGcusjrahG5sZ/fG
AkVGGp5n2nctCp6tF1MldLNJHjzc9smtYt4g/KNil7zzbs7r+EXrMEKx1aIavtfH
icvsqvOniZn8EnkSPj+K/k4aPVjSBxJW0AwH7YuHdPaGNYhc/HDstYKXfs8cD5cY
f2Tm1gzaVBNBsn4EWQrKfUw3OOHACfAk2FwwuW5sCuuVfWASNQ3VXd5hqlewZbk4
jQt2J+itnhCcWZvqN81RhKP1mUkm4IASzmCsyDVyLpMG6hbrdA6FZ7YRfjYR+Obf
Lfcc0g605pxCVGtWIKixJn+A2W+JluxbwsOqPVyM7XrmsHLLK6LOGK3voerpcTwo
tZUJQYuUQVli9edmHerGpsvzCINKp1PspZPPtcqjotIOvSsJ6hNKXDX3CCfQ86Yx
Y5n3GRKiHKcJek/ZAtfc7MumSO+rqd6fO9QwI4MqixBjkOcDYsuKmcdfjMFWpfDF
6z0dmCSk1zoquITrWHmbFjR1RHu3EzrP6lQsD7tVENBKnOI/+LBxNhxsCOwsbwVe
BfLeb0iaii32rAYMDvTHAvrYAywMjtU63wn+seaYIaNjjzsKpoe/RByAYibLg6lN
Ha0GIeK+j0QV9oPTc60LVhy+nSEiZJSCIK7CiEotiR3JJ1ZgdcR4ioAMMzgSyRH0
CyZrKZpwrI25ls3y6cNLrCa0mxmAiSVnAuHkgeM8e16uaPHKGbACpkWzWBelvm0R
o9Ev+yfn0VZSFR5yBpkVViBK6EAbOt+Xb5b4HsP2whCD5sL0hPeAuTNOKdf3IXK3
IkM3ItJIA1nQTwoeMkeP0Y7sBJ7DVtZgxWh09tHF7MznpvFEVfjcM82DwYEIR7ph
/GsOvWxbNRDf5DHv+Uk5VfpsOjP/Etl25+aHUOR17GDbtbWXli6e9UAfPRvIAe7V
qHNlmtqmbLFxHkDEYBP8dVMC/7gi1rjD9GJyTZ583R6YiPu7VaZGJf0guveFwcRO
uHhz+sXGyX4J+YDXzjLDY6n1qQrYiLC2Z7GemWsO2/CXHDk3gxb3UZ1mSktW/kTZ
F4YG9h2Dif+0nGgMKiARJ6Av8kVyEB7hgl9pej8zcpmBm7IIGAL25Vi8LgEhV4ik
yQm5lfgkMTqsg8jwZZYsYjkaQqFsXVlgHGOtacBnkkShL9AM5MGIzdhae0g2uaWf
dR/Csu42elL0ja2ZfY21m+ectIpRpg/H9v2tuFZUITdFuKVa5LXMzRaGfdNUu7oA
ZGUtTo0zyhFiVfDPjUWJIg6MdTLJSXkAUkL7jRP2LxA/FGnnWIkJsaRV5iMJA+9X
1V9OkDS97inJJoYD125oX4m45a6216L0opxCFDnY+yySdh/4bATxM96vQquWfAkz
oICeIESLa/n0dg8J4NGgeQXE0ven9YvNr2IA8ZAgm80bTKFJJrMtyEHBlFPe9xuV
rg7kWdkJHo2Q6zYRKXPgsglbMfv8cfGGvMex0l+AbTkVQfkGAj91DXJz6EsB+ktA
M1smOJkpbK69jBaJPnfZbBzG7D0+/gA1W8uczNUnuZm6uzOqyZmvgRwTYS88PHB7
+7czGT1Q6uCWoRxtJ7SVvevaubNNpLlsT1MmDRzV0lGNg6RVARAeDCBI8ZoHZN8o
0azAFK4OxL5p9PVy9VhyCwGtducV0sfbqh7WICtcCnkv2vBi0xyENzG5cFqLe6H9
QPAU4PKrRN+K+m+PsCAu3bKGXCHSx8R4SJ4iv1rxQeXZRa2p9gSbFrTYkaN/Ev15
Jt7mZoIcU6V5Acx1AgVW0z/M1OwktQZBK77hYXAp7N0Wiquf1YH1MoA6CDIucNvp
zi9h0585gmsu4QrSXbreQBT2LVhrzkoiOfsp01taxCoGHtGlt+donNo/EU7m6vJl
0+V2Gml/9kZIKzJAKcNzp7K66fk+bP5i3qwvVoRodf+fDzIXx/xOIdICcGHVuQW1
rRVU3xCHKhpRK/l6ijufxyfLjOLCSjkvFir5QrieplY5m3YrtlxMs9hqHr8sO3Ir
VEQnXeSUgpbV0DdtPRX7GmcD0VFB2i2UjtkCiXCeJgdpI+fDakvN/e2zLZeXFzkf
Oo1TNApxkh6GRY7JlHqNoErRi+HLZcwv8pD+rrTc9W+5BJYpcttDXatmuLiOnSSR
FLbVnljsUIcogcZHwm6ZS9jpskCcA+RoUA8bkJcGS9LHiGJ6IJNhgwQYjlQfhGNM
aDNu4NmOgs0NQdTmToUSL8q7kx3P4uYh0AD/C5hDQEQvC3/GLUBMc+fYB3MgreUw
Oj/jRoLrXhVdvDLmw/bn5ceyAfOFe+K/Oz7q/CQUfIRzGOpsjXC8gbk79C/fDo9/
IILjSo8+6yO8BgzcwrosLgunfUBM6CVneMbZdCt+j9Ha5Hl28FL4xRwXKPemDzDD
nbc5KFWu3rOvF9IhYiiAtUbxRbhKGsteQPNbsJ9buUpwBvzdoKhRKhxab7jfyc/K
h5vbcRlTIkVBFoIOv9UyB1LmMtY94sSNt+IS5sf1I0eqq0mXBWY7yh17iZDOJOk2
fv4UPZC+6FKUV9h/WaLdkdVHZE0uP9ml0tdLMRQULiGdNdJselEDMZkucMdjNIvr
VkWNInQ68S1s6VVqzEFYpZamd5LdtaNU/c2u/tHUrg1Sb3TJsO5IudXV1xHlhLbN
D97ptPbfdBA9ZJjMWyRMseokWdEkLAzUcCiPCAMq+fT6NwvcXmAD18HELdWieUWa
ouaY+uWv8vzwLVerOOKURBbONQTnjE+o7bEvF+tzIa8UbVUdzudGncvQQAq9KOiD
dXWF8aj1xTYehUZnoOG7Tw9pftAUr0xJ3z+nYmYAUeX6mGteZ8Xm4PJe7w3m343Q
MN/BbXmqUqARCvitjw0MbdtZaukXyNNpiNy8bO2Muuzd287S2KVnvmEHnwFumnf0
S9pkvwk/JdjmE7p5ahftt8i4RJGQAN4l7PpwDNPk48Cu8yhMVru8B+qDGHooAOoT
F0oyY1AIjIxZJc4epot1iLKBAAbGwQoUggN15gWVha+4Di0sUg/pbTQ4tkqpi9Rh
K5uf8bt25oPTfRAlIg6QdvyRc4mm44rCsb12DMjFHXsNG9axUHuOUr5l9mdsuNTS
1LkXr7oYe6HrKH+XR+ky0hHZGKCOSXtnQrUgHQv1hQ1BDEBARF8QWnyYA8Me1qY/
oRpqwFY3SGyjrEVE8hVoHZJqlVXb14xzeJzYRviwMuFfoenP+CX/bIEv2ibPg9jr
FlvM6Cywmz5goeWho6CmCEWxaCN2EWUV87MvrxA3W3F/VOJbh2vLgPYL/CnTvv7V
2TOYhoQFy1QM2yJp1BgULrUmmy+lY4MzjQWq+lsTRk3yBcbQwmuadZHTf90vEUKQ
XApKjystb8QJjtzMTlmaX53ELSO5xCuyTmhry9mvBAqXDZYqRz8Wmya9RksLGZWT
2nihS7GiDTGMTqYKJEjE7Ycv7Sxp/wsguw7NbfcIzYSspQGMaRJwojBSSuYoe17R
P70kX36qQfMfBE+uj5tC8Cnkq09ZzHqdvQzPXaf/bTupr4U2vPMjbWtgUPjYOHqg
+C481KM4nzfFVU5oi0NIHQw5tBJC3RhJk2AxdxDNa/2htwo3yyVb+hqGz8qg+NTF
kh+vG47wuuoFIe1GhSg2Jwkw2z1ZjjiCKQxfn1yk5mBnx9ZmHEWOJQ06XBvs3ZED
OgjMOOEq7LYXO3I4g/nQ2TBMe2Nzbf5tSEXZv1++8qUysNH2AevSEZ6q+DSSg7yB
tjow+05rN1eh50bmMg0iDtbIiPlgspaBlKjSiX0popWuHKljMrPbptCoQdQAM6X+
wS8yMbpvEs3v04Fg5t7wN5ulBbtuMhcw6SxN57iK4ysfqDH5q2BFs9Xqop25msOU
Pj6DodtPVtW3iT4geGRW8PKrDMNGtgc4K7IdI6rA3hsCWPIGVXPpVi5wFQ94Tb7C
GmE1biybcsG2w/cd1zA3hJ5mHV+1UIqKudpAWBQCR3HU60kEPbLijSrFahyDfo1D
44HWfZ2LNunfRCCcbxOaM3vRd1wAlLSiEJ5/wMj+8ZC7OpKhHamnUMmEqA4O8Nuo
rO2gecAPlvfbNmsrkgnNiVtDhuDFWN0KE4YgRFi+kFWMAx4rQ92zhHeqalUNV0Be
nrEEE4RdLo68IbvIXDQaveaEUihcT84vNxaz2fRF0Hv2sml8YTDLuUVkU5KEjfB4
PJHSu3WlAFHch7AgU0jhS0VUAQ53ndh8tb/GkFdd/CFQkwkFwOYBCXA+FYDKDZRs
HPNKq2OGRY35rMhqcpGU0GW+aH87iCe07j0S0yw7IHPdoborFhduGy1qmNJqIcsC
PH1GuS82eGj/cmEAWM9VbIZkJOWQkvMsCnj8WTR4U6EktChYydkdvusU5F6aWj15
Ufu3H4G8egspVhGXNv4X9xBsiHPg2/7G+10OFFsrRndbol4ypfGLAnagvffduWB4
xTMMJ7bZ/1wEgz5NcWXAggW40+XP3jwtgXy4DbjabKGuu9rxhoqsS8ARM/JhX7rj
8mZ2poesRgShWGeXBabCjwQP+Jtge68YcXD8RYDTo9co1UwEwhgpMv2dhb9Zp384
rD2lOqI4//llC3/sUTc2OQAqOfAAen8iGedw/7uu0nFoJpG8XudbWJWv0rcerRzl
hYWe2mTokb1oj6IDvfy394L5XktVJiYqeozsmT+kQEeALo+3SqHe4345VoPQ9NTL
9ebvJfNVwGE2D8htVFuvL3Pt5uR9ZEeQlJ6NUueHb1u/LvLwEHeZ2fbq894j+Uwk
BopPtnfaOqaw4d9i0XWgYyyXHVAWqWMWw8lmOBwCIjtPwIXd6gLOv4o+cR18mxl+
RrCV79UjXPK1PbYoOgLoOcVQSsrd3VO+UM2DPI6A/Ni9HH53X2rf5f61QFoOQ0MO
N0nhw6+vKnB/vjaEtAG0AIyhxbt1N/7UoZo8JxJuW2SkHppf5rWM0L2lyt+m4dnF
nh/eq0nDj70/jrDkDHiGj0qVBHI9by4GFbVzr0nvDE9ad901SnVVDz7ChgL+geZS
EaPM1MJby6HIdFf8EpQiHvZnzQTmDlAUV2/Ge/B3bxX3Iu5oJEoQ6H+1s9fs597+
GIkZAGPGptMLdkmJPnhkLUBCljiHpBseWY7lMGryCsNedbIBfzxg+fwmMx+dhNP2
ALIpmJgrrI160SVq1Aog3AstQP88tPF8wNt7GrtAXMD7D0LQnUh13+G/cx8gi4MD
M20hO50RK4Rin1NsmDabbPnVUxAulh+ZmpVhiARR8ecN1Ux2q2n30V/cVzfmu2E5
p7BI8pyJHexGLxwMTLezVrAYwVEGVzJNp94Gz+nuQ7aRhgiUqXFU/Lm+trNbUBbk
Y5WO3BkGpEbPOUb5XhevgKcRCqYG/jOLDmro5OoF3DZccXkoyrSdG86uBzpuYGAy
arv1b6hv6AfgNZk3fLyAy9pXgTfAiDYmQYeouHCUhpfNMRA/xrYs/YnmWGmNwq15
ruT9BvGTOvKews/kzwBH2k/92J8JauAJyUOhK6Dl1ky6qX1POLqcnmS9O1RFlZ2G
it+afmfwqz+bSxhfPFr648qazmL0J/7iJ37oERBFq5M3+l/WMrIE+p8sy5N8PwPx
jG3jY5rhuYSyNXjxG+RbSa2CaZhcDSHUPooVUBzNbcvuUhxHZEul51bkRKTT2lkL
xWkL6a7Uc4RCDt962hvozfEoPvpCPhbUhwiCXoK/qtzKqvkQSH5UAl5VN0H7MLq5
chHUteMkh9kvL40O/8ktxaD/YDUPpkaIuPp9RCSrBkeyocjcqcW73t0WSbQCyvzu
YS85mUkY347eqxr1omYDs2SRryWNOGHPkWQTLZKvSaUtasO2fZIohTq2UK3+EXVn
xm0kHGEifAPhSph7I6cyCkgMNk4pqe06C21vdm86AvJbYN1u4KPiSwVmcVmOBptP
mK9lx4pcZe+cQDxrjUp8AupHGbKwVBMaa9uD2AfPk+ew3WxvE7X2CceYK7jMEXDj
jWP1L07C+fcf74xKs5yj+2OvL3ollZq7TQAo1hIpQ8VInsqtQniYXltMKXMnWqT6
8cy9lW4K5lbsbmSJwKRBsisX0UPDn6lUrBRRAvq1KFmNlj0K+1HpAtWrdl7x/A8x
rMYSwy0UU/4O2kZvGLl+Mo8gdB+KGpenkTg7LOYa/GKxL/LWvBkl1l6cNhr4rKKI
XOegD6ZONFHJYc5kHBAV6zXhQIWzoVH44aO8gHOCkULIN40k/wJCb0iYZT8r+uzR
ZGtXkaHBr4m0RO2SaLxnhK67ExaXr04iCxQmCq0IZu42y8/9aIGIw9TynkVHCPu4
TtGb6HwF8Fbqe0gbdNdwJVkIQ0NA42zSKBHMaFwmZd3EJDR2exrLnTgN+vWcRC/j
G8MuTADPEYnb6k7jHeAAnVkDrjYTUarnIrLzpCJIpzVnphryinHD/ca1TaLMrAFd
ETqnDim53nVcAr/LJmFpWLBrEzVo5IPYpTihqmpE2BHDm2ej7X+pokCHH45ideK6
kFe6h6d50g9/TiKbD1NvXNjk8oOt3NmI7hxQ5ILe6OgYOKicLGK7zWPO6MymII/r
qresqkELPG4MJSymB6MJ+fshlBQKj8wp66t/4WmACHmLgsB9gpCTX1G4H5AbGWA7
r+lbqFKVdGgTPk8DtCaoit9TbA6kZFRBe+8NfKeKgAWs6+XoCWdUZ8GO3NeefPHS
4nhyHo1xUr8nseJp2chBVnGz/Mf2k/HCnBlKY17Yb+lZs87DyAKQANGEDfgyyFP3
zJtAWJJiQ7PQT8gguwR2/NwJw5nFTnIGrNBSuhY+HcKsSqGbj9/GtbMcbhg+jWBb
AVqQSwBkIw5yoYXYhGivmFjH4jsH1aNPlDp3V/F/tS+EAlQTSNrI6VG3aqnmawAY
JOO5f1Exp2Ucpjue8YMYZfuKzu1mihmfMd/TXf+G46FU5T0D8F8mp7hhrvHWYL2J
Liy0u02uHJNrhoDz5orPJ8IKKjS5m0rz4csGFhxHVX7phisIL45nPf8ZhlogteEA
ckiGekEwqGjCi38In+SRdH83qWfXmqujG5VdxD3q/Tab83E2gSQrzo1/hBLUUh+7
nxb7xixOa0QYnXNoE7SYvXC1lLLZX8zWEcGxm9YuMAjweEeNQlTDu52u9K4BVmyZ
5BfwSnV5+Z3H32JcNTvifNfj89fidEIH2EEg0LomABXgA0vb5TImSRthX84LNd5W
tzoriqgTgfJ7sHoyoAijcYRbcLQuWOxQVJXlvt+i4cyxfNxy26vvg2A/fvsZFa3T
38nqtO2ewZr9O6jdxRaWHLJjHhPsGBKmrSBTPgTp0mu9Dt1c/3olcfWTOHiJMP1Q
gEhX8cWjMLHTf+G3iXCWYcu455DcFdlaQg/DW9jj1sAJYP1oK5NiF3ySrGX7HFQS
8cU61F9M9ezVOT1kvzbRqUVu/bQ83F19up6QKt5tpfLNB/WmElFNRQbRgXFvyxDp
DOAB6sTj0fXyylC3udSxAyg+4kuQTJ6xeOE+ReOY/sLhwiOeqodKBnWrd8A/Ayt1
f6PHEf+hpumhqaTb15uqvs+vb3+5wKwcQa9A4zA5XqU6wOA9XMTWkojH0N4SUcuG
9OKvWrWMAJryo8Gmvsyb4+pYMV+WN5vE3LGFFSWrv/MfHe5HGaGhkomq9p3udKhT
LqptL1d4+xSk1QAqEBGYefk2zuVZPOxMurkJ/lgUZTvVrSvaXZBdbpqTF5Skiz7O
vWL9gjyNkahIk4PRZxLJQozYNitJPdZMgXduazSQ06Rrl3XE0laTQ2AELygNuPC1
Ben4F/MeafLvWl58LTrFLpenh7fsahOoJhiolieBINYQre0PMEeIv9/xUzb3A1ja
mxPVUz2CYrs7XuiHlw2EY54Zp4jajqwZ5bKDUuLRldD3Vh5w5emTPtF+pPilCjya
w2FM/ve4GvkwK2i4I/dwBcRRCCwA2l7pkT7Y3lMEWWZlrZBU7b74SVwOIaiZs2H0
3R9s0alD1tkSTQ14bWYZyF6A/WshjJFptbVXfr6VfnziC0AZwbrb9FAY3uRhTA+4
m4n00eaE09xHRrUEMduM3/2xMTrzcW4Mt++i7LpJGXjkzhqNhtlBQsj2gCT8pNcc
2l7DcT1JigWKT5desVGFUhlbWE98CQT6VglHVRKvwbxbGrYYKe5GNYepxE1UidBA
BteyJYkYi/D3LULMxdZ2h4LxSL1CBm/PA8juqum6NDtDoXuUfLvgNKBc1IdNl1aY
SHo1gB/SE4F3+EsrgNGaC2T40lirD0bQedqLheeibJ+t4Lcmc6UudN2reBWdQd7S
umkt/fdxX2qSszK4XnMVVmKA2KMsKrxNCyCtTyCOS3aMFBMK+Q1l34+P6fELELBM
R3B/f9HccjLwjEzKRmAGMT9+97yeKk+Bqcehbnj2dBkR8TmAO657tkU02wSBpQC1
HSoTJYUHwN2XM75fcpcAIZ0NwUJwyITu0D9I/sXg7qD2pETvxTZcn7tSz23WZTCp
ZgJk8oAVnPJQDSeLIObe9ohh74pIj6cno43y7KuVLDkPLAUw2tasWMtjYPRNF4Qz
/DuDCkfGV2y908/BfNfGKGTjVV8L0Qa5t75juppWD6dUfAGCNR7kIe5Xa2fk5Kcg
fT24tOTYDswANZwIYTy3j6hDFfbUEvY78JyxcBZHxOySxJhMWNgq8qBO7/74XXb3
AM5CvFhaRNvl6JCcMDVrIWE1D3L0ADQCmuhCTbHG4yggM4BY9Oisid4lRMBvJFqB
guRMUcHkvgrxQ40ixbCjnO4n2z6ci/jbsmX/MvcKcWxuLE6x33JJYOV8Yz+icTq7
1NvRxJ4qWIQgqdnLlUlxyP9pMuoOrJspWC21sb0yXmUTd44qtd29F23rlvySTbax
eWCYnOSrMtCEnwmSuWqhvrxFgyXRa8silUPAqimxFU1yNgwa0UjQmT2JkNfyz8hi
KWOYJSNQje3cBstzj1wtGfiJ9lYTAfSL3DoiNokvTi4EUGhxUzhVWT1L+9xAcKAd
mOOfEaklAye4+CJJOWoNO8P1OK3SYvlEVImcmB/kQ1V6ay8byf7HUcug3qAlGhFF
YBC8Hgz4Bg8c3Ui8L/iYVR3bhI/mWZBfzNHWfh0Q+K43k9Zc7pESQG9XXGtb0Uv6
U6/G6Tqf2Ums0bvaNc2aP0/GClfrtOgWFMZpxbOdl/geIZu+JXa1AeLrPZtMjE2x
d4ENFZFuo160Ogus7yH0qWi80RsCRezivii3z+RBpwBkp7OAWlVGsMg+bY7TVAyD
0TFM17EAOHEXWbcXKAWQ7dIBKQKNHOfoKUMt5mnR74NO6Jz2Oqas3IJaUDyl3x3C
eNWFeNaUU8e+mGNcdwx8x+9Ig/ZB5mPWnrmXUJK3X53UMmHfNZCnGh6dtRhjbNXx
MJ5bdBrslXeVBBwY9Q4+64XvIPfyRmT3/nkBp14+mTH+wPp6BIjHCexMw5XuOrD4
NnY0y1LbutA/mEiO9uWMh+ct1su4kPIYFDOFKCJKypIz/0IIi+9C6ytqxMnV4gfJ
5FJ3Wn9yE8xjgoBJAe7vq62j5Xq8wbh6GF4rZVyCDFLMVP+Fpb1A0P9/c15M9wsi
qH02s36vhrrfDeTMxEfxjQ3OTNN2VnJTMjgNwsycINnI8XBRcDXi1wrMn7PXDTrj
acKNnWF7Wa2rascOEePSYa5x9shcVMhyBPQRi8hXSzwXrrBOZS/LKIjC91RoIbK3
YOvZiJCVNMn4WeOMIxidKvq5XJFkeXSErUiP0FpvtsgFN3GkIU1F396w3paiWMEZ
RuGROuQFB204e9LnJJ2K2XVPJ2ZlTS7EC5N6QAK8IhnIvFkyoAIJ/F9x5WyvH5Sy
NgvTVNBPEDgpGKZThuFlUdPih4ejXiIXJBhyGQMj/qRP3Sv6CY99lfnhrLdFuisO
w+lP5QhhJwq453r3iKSNrXqKpWEl3kyTc53SS3lOm68r7QmGO5s8Sp1TzAG1jn8g
D44rKWNX+rWlL4aKhqYk0i27WKeQ11SOzpJt37B/Et/BFMGQWbcJb8m2ApSs3FEI
a1hWJVY5MtS1twhV7ptVlHTma2JQFsRVh1VtoEmzsWl8Np1oUC0np2F5JIhkIEfn
0fOSptpM18IEVbBZNM/vpGrnMrsAAmgOFei7+slWftxlpvLA75eoFV5y3aZ7e6hg
3LA9x+DlJY1MKQx45er0cbZuDVtcIPiCT06fGlBrU8Xi6MNgLqdzA0JnFnDf/Rov
pyX6MLQJCPjqaABreJfR62jwPf3E3w2rLGT34yjtw/WsnYpJXRYm/Yv1O/UY+ZYO
eXRNihisZ+gRrwpNZe863HxWR7sP7hM7iVi1lVZNU2+ARhDnGCMFuZwlCENrzp0l
lNYCU/phIFWBjOPeKXWXPk5uUKXtQGqJ88O+2lLMulgLi6RDBcgFjhJGKGCTREdy
DE7ad1wuWmmqyCPWg7JNlIASflXRDUn4eha2YriSiTY14HsMq2ZVXLQUFocsFObL
vRTWNLZHmpbx8FPn3OCbJZYjV0CXk4Y2d3BvvYRdKitbnmhpqo5dtIoVak/CAt2N
VYZGjcdEQ4sv14CpSzlOoK6MHMjk8q8/nylby+O2BhRrNgmS8jNK8MPWGc6Xdc2+
kASN8UZIIdOOEvG/Wy2F+4QAtWm6OOxesMjOvTc/nB00HnNVmje8oZiQR6uaaCf0
SfJvCbs5gPXFKJm3sdh8eVLZF6XMSqFAwAVFVJSw/xQ6EZvQg5cyoctIbODki2PZ
gpmQlaGK578OFRTKY6kiQ9vtMhJXuX7CgqWOrpgs/mpzRRpHvcJCFJ2EBBH0wFJY
PyxiUhjvZsPlvc/SROney+PCG+SVoND2G9V3teoWAULljeLeSzwRj9JSqkTVnFg0
egf8Bhz6hkRi/d76LZ7bNSqlwhnGrDSVX7XXcOHmXsUluLRc/3bkJFpmaJsXvNfn
dFa5hsfal5hxfgOk7R+Xj/CxiNYsjMb0k0dnTEz7XEyYTE+fFBUekaIeqhZwi1TY
qevECEzAwZTa9QE1wm8CUxUHNuCh/jWVadjL4JN1vE0O36Obb/sehGr05eZ5hkCn
ilrjFJw6NU/0APqt9t+/85eehA/UcFVCknULumQ+ONJST3OSQnu8h17drwxB7M9i
YS9V4CQggmbgr3rX0BBLX7bh8AIRIg8MbXIuCAuqbYo8h9LDPnlCNyKEV1No6BRD
F2Q0yzO34KBSckhhSqA0FOfF701JO4WYFCT4b3xgfg1HJsaOQ0rtRVUmfJDPCU5J
NzyLHWLqKp1uLx5/wguk7bwIQN8WviyVoslqSreQN+4+XS62TBE7aB24jc/b+pee
Wm81fqQt/C685BL0fR2FjX+EG3ZoWLMBJuNIiVQwPa5eCf2dXQacdDrF+v90sKqP
DgWSYdOdMEuNwxnzqEOxAFyVgOZXdne6DHFVuKlIU+RQOhbdrfHIQtBACWcMz5RQ
9t2QSemGAcr6OuwW/HT4peNwAUX6HoLIYJYemUWGW0F85Fsv9qf6ehfWa0RZaoWB
8qVNCsX+zxUie2A5c9ppzgXyArsV4HgqUYmWBEVIloWW8px5Wa1fGcKsPUzvzKNK
+pUMyVrJOV8CQrx4YZWq2BLqylJ0y9tJZOA6OvbyS6JofvGQ/4/5iEXnngTE2Ny9
awt45kga0Mi5wHVZTXhO4MFo2AdzKPfopgH23bvp2CL7aFYFObojQ3+hZjH3p+Yt
3QU83Jii5h+3olzGt4leHKYRB/GJuqMhHygepsKOjACN29RavU+tHuzBartysJwo
SNuZzI6Ba+uMKjorCVHqwfPLz5buFnBWYr/W8DRrGABhdsOHpr614tYjanwDrzdP
sqcrDUwic0vZGJYhq61kcb7rYSypdYzQ6w65XWqGFZDMrK4Zzq+G7PbVYKJTUHNe
FOZ3GSKoR/u9Rqw8k8NzpNuGO7pG8Fj8qxj87HPi8rHbVZgcabu5MgjE58PkMkVe
fu8gGPNyH+97naiXV/SfULw4tc8/8By0u+9tI3l5lF7wyjsk2pn85X0TAWmMRfwv
R7O5DV0yORHGWRzIcZMNHMvCD+IN9NLDaCWxWE7B63+cUEBJp5VoEdzEC0lHl+cr
h9uLtYOMmfObj4WN5X50XK0WQKZSRidJVg8of+NCABPTWswZP+v/+cDnSKXCr0zS
+QmsrbBWvLyvOf35s3KbEtvNzQKMZ+fFfXGrcEXHxGZ54PvQWEgvZIVKIV+hPxNI
KCZzh9lLHsSrOCuS1z3aBGYefpxbl1z5MP+FgfMN/wUzxgMAIvqG5qWjhNsU4Ko+
J3ntO0QOCqzsVmywZwlQxUrKzaexiZw+6dHSPao7omHmgvplWqpfvDIqdU/rF2We
nEdz9aNPsbIvibyGdl9TNSx/mbXwfGc0DQJHCFz3md1TMQ87fpEHyZlxH2xkJNWX
o5gbW7jF1e7Z7Ux92OCqVli2BwTXEGN5ExHryA8+X7THq4h/gInxu+7Mo0ag4Xuy
I4gHqYbdyo8tIKLMMF+Bu0XRp/wV5Qs/9SVW5OPMVxV/+joeUDxvlCv9PmKKrczC
KtLDtZD02UNfgKamWH3+Ne6ABn+LIzw01x2Gk9AaWTdW6rG1eGFW91ocolkNKFKK
LPHogCA14qxgghEuQbCn+11wX355IFKKzyyPejFW633cpxkz+/3+zFL2AXnpkDPn
OBp3ts28Gy9LWyMmpjm6c3XZyHG0TGzjsnVqcjGQbqPVNohmYu5+Afl7GMDXzZqS
DyiPtDy+e3W5m/mR9ozY13+/z07xcnrJSew3EZiN6EDjBe7XkdB0e5A3V+8vE/aS
VkK0TPF2Q6z+zq6jThuN4Mr5iGHrNAxqOhjEAokjev65RF8FJQy51gk9Jkvm3sJw
PXoO8k0AdQdUWt14z78g/P2uP++mMILXOagC/B0tre5UBWXlMfHRbof6hhW4hvG1
kEH5QpDaqti+wAu7PPfMAlVehfM65GVG8WhiS19NgjE6tQvg/FW2Eaf/iQMiXC7/
uf3GgaIITo5sC9NC6t7n26jg1l1+kSycK7LUGN5+XQfmtzCZtDr+bzpbHi1j0Gcu
9IKo9BTxttKpDVX8a3NuK+41n1A4Z4PSidAlTZgVm53Cjl6aeQxvudbxGkAQRir2
koAUKuZnWb8THdhBNQJhkgfr4ZWhF49CaJcRJoi/cKgKTC+xD10AwgigqcVT2IXb
RAFTFZ2kW5c4TVUBvWey4ChIiOzeU6BvLmrb/U2bgtc1WOyoTec8v0R8OBS1GHLJ
3G1qDnNNNUIgK3eNtvc6jNEkSn5e1WwcOdMLqFZZnWfuBmQvk8CAfrXJII6AWOzO
NYXw3XFCVxbpRhE61xWbqI9uWs+DGMoFCShX3kFXwjvg8FNaapt0oxdIJjXDlpgT
TfTBdtM2hvT3vJoOnbJ3uwtVHp4JFI/Hm58G/vLyu1QGk2mS18QLn8wVU7eS54rP
Uc75IIjpLpF9GYsR2FW8z44Mc7E5ihRxQakG1AckcVIWaOZpyx0lr6Lhx/2lyNC9
k/07NLaUSndZB29yh31t0c/VFyb7Zz/CcQPXNnexlN0boYAZa8o01TpxvJFd8A5h
g2rgVJmyqqMKqAn/4pONO1bV+5D6x50k8r0IiHzRpnavapQJj67lHprx8yyeAPKQ
0uQMdDjyl6A3n2g6B6wkdyt8CHHa5+2o6k2Jv9iwsHfILxziV/bpQEH4TvsCGz0J
tKBvcorS2elxN/PwIPkpCGpefF+gjo3Jmg8MhatfzDgzRLtBxpxEbS9ihtckdCst
p9JN+DFhllCLzr1f94ZGHFmyF13iQjkaGxkNMb+o76FkB71WjsG+OCWINzcx7g/A
UoCNU5k4aTwVzobBaUEvfue6GlZWg0fo8edmqn0N1MbSPP7fmuSoZ7Eza2ye9ziK
fK0mWYwxuXcKSKd/ZlN6+ZKzpv29HsRDYr+JTr67L+KJ2HAuwwE78QWsKeM0V3rr
iFPB8Fx/dlShizNpSXFzJE4VReuHf22nRlKNIPjFFdyr3OPs9yY8kVJjSgpO0Lcd
M6ooRSiRITKj9v+waIizW/ICrAoekDQpoV2gjZpfusa5WB+hr9l8p5F+ePBOkm+8
hAXe/c7HZL9kGoICCnWUPp0TC6rCR76UrLJD3P+C+7I/P7mDOZtS44OsrEmdo8X+
iRMvDAUlJMH+KWta7lymr1UI5xTUFXKWirYpwf+YeTMXzUi/s6Te1xZcJgJHEnRS
Oa4r4R240tiRMUlhUmdhvXLnqZHY3fcyJqFPj0iE9X/R1dOO9LkNyY+TnPNlON7p
msDQtnubAWLCVtxKxMBUlDEkRN5UyglA4RXEWi0wSW4BngIZuLV1TXUXylywACJq
xV4BFGcYxZlhIDqsU+snnSGzuOrX9kkKlOKuA+eFh9uSJDyLVQ6EMOwly7hBSQBM
udZdlf9hntbGukE45ZdKx29AlqrKOZoICfeRS9C7r4UGXQGg2bbNvpcujLnSL6bJ
qBMvwyLyhRIyeEoYe7XcoaoH2GVR1K5ubA1AWE16JRCd71YqDbg2BCt68lg+inSZ
BuF7a5bHifpv94Q0l1dBMVedQE1+O7m4hx9zecQTFuLbiyERI3MdFXKPx1fzO5bR
Bbz3LSDn9bYy9s/na6+1TOxGCiufZD0zfyJC87ESuIi+6r2J5OBqITHzDVskmW9c
Bj/B/rVjNKsXivxQeKfp7ml0kvUQg5dn7d8moVqUW5HYJXPdkK6csUx8tF6FImU8
CC008twAPixErx+YhB+xPa2QbJLkYsS1NTw/HO16+OZ+5Kr1b6L7QTCHoLOsslQM
xC8Iuws38wtQGVCaqP1BwcjS8nHrr/HF3Xaj40/tuLgrzV0qZkXMcA2bEO9WIZBj
FPZiiKJQbg8YrrNL/Mejfmxno/TDjs8eZnuXyEuBsyaeawnmybSUK/kU1iawgR5u
t0eG2cij3+rUj+FT6TiNTHHzgoscR+ipDso7tToYf+NNrR2geaybL9Tx9q6T9JvJ
3Bg74IUUDErkLXd96zGzustuhZNoxFomEyw/5tDtZRkKi6lwXIO9gquf/APxUcLZ
GPjktrEgRaAm1XkjYYowotALIyJo3xnVMNKt4Degfyc20v8U+o/KKgjbgnrY/AHv
V3VbigwXerlbJhvuJj06vV2N7jmQ4oy3NbJTjqnmlDKty5f4lXyvJuQbtik1EgsW
VaZaUrQGL52jtanIs7w1bdUY3d8G606vp6szSTHRI8EOJlUx3flHadD9Znr5Q01f
D6i0Lvdf0TEd9xyU7yMHqqA4a4fLx9iKT5h/ESDdmNi9vJAmZrTPdZApP/MrpbTE
sGLten2MFJcYfkOqbaOkquLuk+yTx61Lq1QgHDOSsfJ9TSCIvOHvX+E3pKYi0aYT
RKKfPwae1ILhM7rP4vbqy0sO6i7jEFRHqVgpb4/QgK7udbFOpzMlpMy6xlnxkFBN
dyu5E4bkzfS3ah/jqCWYjyQAmU4D3RJtBRnQHSBMsP/zueP16E51JABjh/is+ptN
LP+BqLP+wlpTZ20lBoeSZOWzZPJksGnLNUkOIAzOv4iQ4FcoUSpjJHYNzAYFe9lK
4Rv9Jlb6KoAbHcp8fMAkWOsEVbEXp3QESCGQx9QBMvFN8rGiTVyx0Uc1rRoVExxY
o1KWncLdvYhGyM8jgBw/Ox79KWEGbvYT3qyTLYT+GA5Yumk7jgpxxFa9lyFehZNE
SUxq8WHcnt7HAH+WqqffR1xo8xcF8WRvbXboGQHwgo99Dmq1EkQ9fzSu+Drr1Dl/
/O8EjcX4WP6tIS4zHU8lnl7Vp4oLUp1en4w1ZDcYwJVOoxPuuqLJJvBMmatBSxeZ
0tXmBgG4VMHGOCDSAXJRlQBJfYiOxEYlImnAHssoe0LgoeDUvW454q4aLf0kS60f
a5Nq880zLmlRk0SwUhBunl+ik53xMuHIJzeEilyfIJjdodIF331E6EDYXkj5+5nJ
cht92r1RNlAMrvptvEQNcKcB7c1qdS/BVk68WH1sNdSFwcMglYU69aHSXzm5CelT
ltp7DzriTOxk3EcV+dnq3/uPzWuYqyfrkTsaRcLBPa8AkGn2+YxWcOiNuDo/5jeo
8XjkILq3lALCsnIIrOGT5gf113s/gBhdZgxvoRzoj2MLFOlfnly9RRL4Lh7Lk1bV
zEkr6NGJRiZz32gATiOjXZjDK5TUoI5dzqlj3Gvu2bmwQ1JScTjjgJ8vnK9/aZfv
orOyx1wJjy7alId8mQpSfSxa4j36XnlzgZcI5gCylOxuNrHrxuZKUhRTj2j3HxMA
xUbARVOXlMxd3nS+VlAA3Kx645II/jv/F7T+gBqRSRGHN7FH3vxSCmo5kbQlR3Nl
IQyDvf6tRygc8PaA0E1GSnpyFQrUe9lowUXuagItoA763pqfbPEre3VMRUpO7jyq
no4LnzpOFq8nWSpR5geGlR784j5BiNfpWz0yROm/6sIzVN+u/D82lAJ85B9l+23w
yuLuMRtprlVkOAkiW+lBj/uWM+FDbX98VDwe63i4Gv3G6oa+jpXTEKwju3S9e+wx
GREpkorDygyWb1qpcrtLcAAgJYiFGBnnR11skIMLbKpJtDOGTfLLArBdkftgYZnr
Z37Yp9A0Mar67DGUQbishjp8n3EE9bUhiycWlW3PhXqE3x4DIsM6XijV19YQEhuY
1GxJRm/J/7wu0OhvsIhobGUw/p3EyHzF25++ytRXNsWrHnKlW4XFenS89OFoKcKL
s5UmW1I+D9tAS+ibXRiysqTZM0RjwAw5zPWHOXqVZKv8U1lih0nzpbasZ/exZvGq
B0jimPrdSfoi5qtrfKgwukMalLy7U6316JazbS87md+xw490NXuePeMkz32VYv1t
h+VJ+3dNLYhc9S8S5EZIA+thJjvSqnspTYDlfYwWF2bZZJm6zTsJCgszlpDZzjQP
WhSSdYy7zL2S3p8DV827k0qfniVQLMtOfnkIqGKmxDmN54cNTAgMKk+9lKruEdlQ
tpd7lXxMx9f0xHlXhhjZ7WQ0Zh8G4ZQNKaG2m82xWT3u6cqHjJGbAbMdBFAzBqBO
YfmbT9WGsZhVzjYgz2h+CdhAmwBb1bEV3hb0liwvwv72zhU42XTFSARb4Ge/i4XM
R5e/bIyDuCEvtwR/1CZF8k6BRIGpeDDKchNcRRiYwsfIaE4dUsZo37zGExVked0B
Ai0ENxjPffYzqE5x6dgsrAJTAk6MjPR6x/eX6uUgydtWNmm73mJgTr1v7uIq1FrR
8wsFmtNc1E/B848yyWauWmVTxGTrh9kfJDqpwx9BabstIDfx0vHtoqVHyh0wDR3O
RCPuC6w34hqUxw1gXWwuuovPvDydmeGC2g6BwKg/JA72aSw8CBUi2C8cJzGhhppz
Etfgc5hmpxKU6i3OuudfupE1fbbAxvooT71yRpe/Y/zpY3vjsKmkIK4cH7K9xRsC
3J6HAiiBj6pbhnxxV+VcprPDk+HO9mEJj4RNdGNsL6gLSRtDnWt/hHjZtFFhr6Ep
VIp5wiXlQ0tsJCMAgpaKlqOkTgCLXIe/eqnerZmE2AADl/MgYOL9j5J5wFD3CMtY
+Z5jOGfGetifPeYMpjROH7owv67+DEBqm9h+alDKT3hHDhusxfbR0SLYfglqdcM6
y//EdIdtOKcadW3Z2DQwgsg2yuhLflmw+jPlRCriceiPGPM7PvEL1aa/coDb1S0+
IvTHwK2O/FxYQULISu9l8TQkmhYn9otGF2v5AVuEVFb7inOLSAYZPnAU6KF2IApp
0GcFhfmVIsTgXRteCFbvI7+rwmj4zbls/wOosabF135fP9sL40gRd6BhJX65WdFk
gQJbig8hlJTTB1eKvPWbASvmfHkCjVM7Fg2m8xzeAcajzBwW+xSMuvOwspFk1Kuv
pnrg9p5wTdCvWmFCQxOHcJNlUC2hgYf7WC+czqzB9Hp91/YT/CFCVrJq9bQSb4si
Zx7X4t8jTdjDA6w6Z8aAORwOh7aE1EFZM5kyKFM7A4XBdMNpCoVqYlwg1kj5BvJu
cEDdQGXJArPXhAJUHZE6MkjH+ygDBQsTNZ6U6oLfuOicZJQZTzYgyZXD/gWG+NJ5
nxQbQLkb/2SBZ2g/c5TpueauVAfvTfs2Sqd4M6lMdUELD+gxHtEAXj9epeR/BR62
VSAo7wPzr1yp6cPA8LhlJBye1FUhdWdgQBjsFgdvsIpQMrtM7GDnVpeOfQCCcH2U
MsM94YP576pXlfmsHxMr14rS6FyRjaGdSnFbVPWDOGed73G7G/DINv13PEwTGlOy
DgUBO2QKyWqLdRtdoQEoEcy1SvGhxVMdQrQuDADcYsLZKm6Fk/ZA20hIemETC+pj
PkVsKyTGWbyzL5opUWXryNuklbkDqHn/yFJ8L8FYc0e9PHJwe6PVYEvak8IqMFbP
PgGFS1+C7oEeOiuT9FzKP4UUf7ktPgxfOf2LQgCD+UR7fDWTYUPiQ7xSZV4Q99rg
l0llQ4NcDlHogVfuY0Q+RflUvyLzSPKDkLcEDc1K2ouemnDJU8n7C221MVBJCfLZ
K2nQ4NNsy+JXp0E4NbV2fhsO3UtEK2NhuOJko0nRLvghx0oGp+mmt056CMMtwRXC
opx3iG4kCu9vV69pP7iJOCf3boEVDxMFRMggrlFbPjmozywzsDZA8KAgDUspbsHR
yoiup5DX5iILp3hvKa4/FarjXp/YSUKE0u5lRrRom4Z9Vz1t6Q9DKKhKw6zmwc2W
+PtK3WYE4dLSkQ0QLojzM2UE4KP+q3yES/Ht55+VFn9syKRa3ePLwYnXkMDp5NaG
DIJRGqqtOEgNVn8a4We9MGUTguNNH25+6xTUp4BHRHhBPmz4SaNkFGK3H4L/ErNP
xzkendOzOAv1KrcTECS9erpOrkHFbWrlSbrEO1TOZY6GzWLG2Xd3AYsob/s2x7TW
Lf9M5gH76y04cD8kVYZRJWayvzJeFrSufiXg9xA0rAgd1xUBuInSlunsmuQyi1gZ
QgocMqifSNlbk7Cm8yWhuKvDb1gdcWjWXC1m1jMqrxQIDRvR3BVzi0a+1XrLE3JE
WN5ezgXc00pnLsre2mqGSSDKBMI67kNxJE99b3SzlWfAtxdZR+gnKPqE4e2wk5gP
eKNJlpNVZaCnmqEJs/pJRrsOzgzBvseYrl+0KtNWPD/OQC1N9k4XTttuSbM5/R9I
oOHKZOUerqAHk5wt11bmaqTXvNzVCJVIzD5qSl/3H2+0MMT2+jgT+sR10zGSEXBJ
Dq9fB/XegkLDIuqGWgROJgO4pl3tA2Ni0Nr7MyS/9KAbb0/ZPR0L8Nu34J6f1v1x
26sPfNr23/r0SYsboMOIl7DUOt6OwdeBOGpQBVrRHYGpYSsffW5cKxrWivgtQKe4
s7YVsEygzkmkgdoc/H9kL3O9b9JX9zP8HGk97C0RDwa/fTII9j++lkw0ePUzXRnR
5y1VAtJdBPUd2WJRw4wmznlguGk94YNbnAAWuLQNA1GnyqOiDGgjBrSCucXdc0N8
Z8wdb40GRmczTp9IfEA5uExuR9aV6COPYxGJTW2H/9XRG77GMcqAZ6Sdqbp792Lu
4zvqmrRCrjOFfQbxyWKWCoyque+DWieLMU3ALPlxktqUPBvQ1YEPMYcnRE01qiza
QT0E3ZJpdPZ9cetiyKr3eJvmxDk2gUSS/PwTIaF9/AJuIOJkjDYA3BsyS0aTTduu
vzuunDDip1VeTFNYAb8z9458wO0OPrV+MIqjKu7aa8kXYALStFFpQK0y9dddWhWo
dCxYYbueVGQjWs+qYoG1LqxsSS9AAksIKuXUZcoOxwGFfRLr3V1FBZDx2eRboKtO
pLnTIkVhSknw1wYPty0Bmz5scgdRMQOQ7HsCw96KMNClS++I1I0mzyVCw/oVeh+G
G7ywLhLJdG6H7YqIw5wpuKmaRIcPR2DHMeDSNfXyM9O1sCm9vHbRGVAcNJVekpuc
ARzsr2LkEGaPyQy81xdXGCUXTLSdLcHrYB5kJVhPdDgsd3pGNP8rBIlBTzHFzm2g
W3/jkUBIFmoynFPbcXaQ7Qd9cw+abT+P9UeJ7CWBXdEkEze8kCC8vZqG0SUbwxbY
dO8KkYr7RITGDfL6DG3RdWnrC/0yQmQJZ8yRU0xU7UKIz3G0d/ynt7A8bL5boExU
lvI0mVJ6dQMbF8mGo4dLzrIDiUktaxniKBCDCgin9pGPUUB0PpOHCKpH88QGChQD
nE88NSNR5kNm6k8lZQWBuP4Ugd5xO26HOXc82kAZoDmVStyXNJwUFKR4LUiHXMAY
Ov7FleQn2xAVaOv4dOgtAafj++kKafJqMPFjWTS/fDsHuue4FUxndKApD0b4oJfC
a/gR1JwpXuINhC37xXai3uymyc1Nxags350ziG2YrNn3sz0gatwW4jrSB6aT9TeU
flEgrBQuq16eZSY2CeL5raK6NUxft11FPSN4N9jFhzUeILjPE5VlXF0on/9BX5oY
fNBiIsV2O2QJavfa/r/0SV8E6CdTmau0xBd0PM/o6Vk5khEy6tVtxbRqZ0QFXdHd
AHmMGTHH8GpblSs0Zgx4C1W3XPhUDlNSgm6vrsCLLx1Gx7McN4OKBsYhf6yboXFm
tfA943QO486lLvy+823NnqOQejoWgMhucPsuKi10A31jA4who3is6tgmFqY0BQjz
tLcaU6/hEAAMnenT5Pg8uLeIIT+J5+ZDKjnVCaJF+QHBKDwFKZ2jqg8Q9J474Zuh
DVZ+TyvFZGdeFUDUdTW00Znftu9v1mxEDO6Z/caBBKayy1QYcO4uqiTr++WC7ZLl
pctN+jGlg4TIHbMpC/LI2KpirRfv5a+wP76z8bB1yXx1bZJfLnyJgrHu+v1xBFGC
E1N0UtZAwhquUl/j+/C2+zweuTYCQJml28gXB5yjF0CUxg6qjwD9Vms5z3s0HIh0
M8nUYpFBvRyP5Zj+yZWmao9A6WG6DMmsQyVMDdJUsQVlyZNt3mM13YdepHQb6ntw
opJozUBVs8KELm1+ExtFdsMQmXS4MmS2BA+l6mOBz9B8Oaw3lQc4Q9ZanHpxNDYO
JCarMOlDGTKG2EXyscuqAkk0I6/h9u6T1wjhaVEvSdNzl12hwarZrwoaw5n5mNaJ
fIsCFCr/sHa8VsBcy78+B50YQ8YOSnch5sD7xvUUSMoqGFQgHnc8Rpf32vDERjrG
jqgRBLxl90MUiqrqlxj580FmGR8BJNnnKkW+ZTCcf1LOIK6qvnBXJ3NvpyzZP5da
GQ8q8h77y8/7hKMcMI/sPVjyHQHe4DDy7RR8pWSJEqby0iVn8KcqudwwnuIL57xb
CZ9/BUt20nJoQi1k4zW9RzNjkNxxJq7cgJ1JIuZC5a+XVXOEmgbEwEu6SMcH45Nt
HNl2s4dNBGjGUsYX8KylbZOtExo4pa34tArjtMTHGn6sRMhK7ERlQuZWgK8520WS
O0Pj8gbS7YWqTaW3Qb2WU5g3pL8j2GgmNhgeETBCdvv/Wxwq+rbXE9YXvIdZcmfS
tV9FkT6v20UjW8UaU2FjS3uZpvaUBEbVfuf3fGmdSeVM2L7EJ7JF2RWrhikgWWhT
3oNR0jFguVKVo15sMh/TqsR6aC39UatRI6olZDL0VaxW6RiTcLsfVtMO7xJc+7LF
0zPHYhFdlSiS++QedQEwYx81NCqlRPD56In1jj8vxBbXuars/kX9MQf/V1vPdNiw
7f7UwY3AT6aqHHIqB51mMk3jEcAko2dZfY/3tpmbnPVfHHjsiSOgVmUPVAHfou1c
qb0/CMtb8d+nDzVajsZc6ixYf+fZXs/qyeAbY1gRFYkcvid3Wm97ylWaRKLSd51x
B1NZqeYQVdwlNcGhpEmd8QXOyjaehALVZR7AfgM6X7SLS8tg411pBDSHoZxNWuiu
s+fW4q1k/kDEBIIwiDLcNuuoKQHwT69A38uDE1E3zvgIG/ny0HNeh0RRpoCEjhzV
psTCc/vO44drfhWvT5SpO0fkDatLPLD/bcXlVRE23uuyi9mQxQxT1uEGuZJibiH4
Rf4s/13C2hggamk6avQmF95e7nBRnkt2EG4bYGcm9z7rDTy6f2y30q2tZtAvXWje
P1g7Q/SNM+uTUMPAtVWofQPTsx/cPS6p1n58d4S/KPk1BVVgvA6B42j1+l/VSHnX
3CEMmI3s9KOPHW4ohMkoBAyPOIIQt3JoXr40+fVSR0cpG9LvB8T/eZDx6dMW0pc4
bKUsGFRm0dtKGjYebPp/Mo57qnl+ha2c00NE0fhMEL0QT69NloUQkM2gIU8RP2SF
vIH8MAhoU8BJvcaEAiLj9HoI/akqw4s8oIambKiStVOQFV7fC5WocFZUdPngPQEb
xL5gAamOvxYs8Jd8hga8febv7k6/zu067GvGUgu+EiC3J975sytGXfrqqBxudIBj
iOa+nivdYsPyqSS0P/Ib4xXUynXkdv/j1iMAsC7kHcUKef6VbR9Pb2ocaXl3Ogcx
FznVqsE44o9ytKjQHVq/5iKdm2L80OaOm1/HcqM71SXpqzoszEopT/vGcpips14/
J4TVkZcswBf3wahabS7x/DMHa/ju/OsaghdnpvL3r5hsXWNwDTKL9DtUCs2nvq4V
l2cHZeZ98JLKsuo8PqHN9jwdTh1G5vXaPpPPofejVxBkOmlYWy3CwlF/OPl5c9dd
9lGA5HlYQi9d8LjzO1FAWYB/n1k/I7QVofXaML7DM/peRml65AB3ToSWLTMzaEqN
UnF3GvmkrGW9LpfsVPDV7KX13cCWQ8bQ7dIvxv/lwXR9WPxWIoHIJFzBzUggwmFx
Ig4MndgR4d69iAxkuTPZd5eqB91dTuykGCK0Tfv05gV5bi9aiBkpisM5rQoX/wWj
7o6BBMW+4FejMbtIyexSxsc8Sd90iWA3BXSPuxXoYv9l1zowvqr4X5kVG9IyGftg
PYrBC/4exB9W66hzUw68vk8JfjCRdM7FGrOZNJoaEAnMBEgIwub2+1kV7X6V+heI
HG8DuAml3bKaRCUOW9ycdPXeXe55iCbvyVzpvFuMBbrF3bwmYpJonLPeZj4pASze
/OSVJuX4a4OMvWqIycUWMfOqL+jj4hs7bDOz5p/O7XBh2bdqfSkU4W9y8EWA8eUS
9SrgdOwergRFXDef6TEpn0Ff2w4ocA0wpvTupUc/soxNBFRoK6oO3Or047+PbjP9
UQbeedKa79K50kyUcVVucYpoj5zYbNGsxLb7BA3qvG/sT9bj4zdGZx3VhzidsgPP
bv63nmcJCdyMEiLIVgi7JnbjpemnIB+4bEuqpBeVcd1tkmsqAARzPapICSIwGLLO
cKhwacwkFctH+rt11QjBYm4jigSZef28vTAf6rYJcAOxQXRbsKJe6JK0gywlAHfr
obMtsrfyKLHlCwd6pfy8WOhbcvt7RAP4Ax9X0hcSDv42vYhkkRFv5ogatJJy8/+S
NQm2qIKXMHd1F8Zp7TN4lWb9MxxpmJwjPcvxwUR9rvN9GTlbi0A39yHlhP4tzvow
Xc7ugTs8iWkfetxDQlawD+Uqb+vcsFfcHbgsYZn1D9mOLzZblWqfwAlva8RN6hY5
qne21gh5440KNRV8ANb5a5+qg2ksWNqNN4Yd9Hyc3kTbPNwU5feOMeK3itKoXbCJ
N4xtD6j+yQdshnfhIimTc8JxUDDCUbYN9bhYhXTv0eBa2SBojq8FtOuKb+s0qVKm
1CkV8wRBCf4clxSGzxTSDq6NiPhkSoTX5tAnMUnrOl0CdexiFBrx4t/03zhs02Lk
SOvyrfe8uKBCSeA1HtlHE0wFLaVtLGVhzt4zwEdoVvpOF1m6T3Cc/mLVCKdcOUfB
Z0eJx5AKZ4nBYxzlfAe08a64TqaccgNgB7Inx4e4P7+nEf7TOE0EcUFSdU2eFYBW
x6CHfZOMJrVDI57ocZ6TDQi8Xpyzr1hK4X2CQwXEpKdkTKOGgFzkhuABrcsAQRbN
iPLUwUGdF58TcxGUcyMNWXHyQBG/ipD6CT3XXzDSKB/1Huft2Hx1pj2bUIfBldz7
bk5yz/gVx+n8qfuWA0O/Gc+Z+w7RIPfdv5J9FaH8iYFsDTnqgJhG1bSE1Pahq0B4
jS8nEEVb9GA/VTVznYUj+fvu4r/D/Uo7h8wrTHEooYRR21y6cSNkH5M2eFYrk/zg
Sm/5Y3FBjeyTYvYNL0K8PLa6BBfWxeU+LSYiwTzRkYLIOTKf0cZvjMAoxaYwvRAv
pRDZeTbNt10Gu8SRbgeXrfKKs9kgx68JNceRev66ImgUYNlfM+s/XqVwlaJX5q80
9aPSEbL9xgssx6JcPodXDkWRToflz+3poryHjgw7bSOGSu0Hn01pA/za+7ksm7LN
3bXss/nDNklYFP4SsZoPCdnNKXqwmPSutQSkuqOR7Edz2UlHSPmb0pDVMssLUHMW
YjZJ3VAoDEouEDmRgvuer8//ey67dZFlX7ogTfALxFaPGz67YRoMVWNIFdoEL0p0
G4PyZqZyEWykVdFZCB0C70TZ/PJPqCmTE0KZHJw1DWKF2B5yuHKCaV2N0euXBjGQ
h4br8c6zxfnIpObhd1pYWfUkUrbEeM2dTzArDgEv8as6ceBpMhHb0aaa53Wi7RaT
YkLr4iHebsiFq3alo8Fy3GjGRM7hZLl/GXQwI/HP6Av/5KGPoZz1bIGUNZesrkAz
yzgqh2UZLPrqV8nevFJIFmBaf7TRBg3VqKnEzTYjmZ9lHkN090XIY8Tk15qD/R+T
dv4osQCT4BEbfw/mOqiN46jKYhR1yX5xUJ1rh6wsg4ekfAxi7m4GnHGuqdVUr2LU
1w9pw9FxzLAs7jA41qTCpif+OnIgBt/JeB9cTaId3bqfg9D85GQ3ocLl3wdxlIKT
qlsURybOSsdlLqE83rdl8V0fgjwDxmJFoInPBO1IhFr9Ki370LYixs/nhR746qcN
9mzR6ZoCQek10WTtKMk32sArg+na7RKHh2HekPiHNgE1g9bJmXz3TgK/8lvCp8Ep
NEv3I4mFk/Vxlr13ce0RVqkNors3P9p84a/vE8gIkIRiRx59QdzjSAqaS77rSlBh
GGiIvzkmawPlo1e/Kh44bF/c4Q5p1ouuWZyMKptYUU1mNcLAm/o5r75jgqhGJJCb
+IIPE7jk5TbrxRnHXX7q1hrhoONpOHl1N0q8CBPfPnsRioNBi05Taq3g2ZcLiIWQ
k0wGnoFrMRBv7MJmdGlw+Zu/FWsYs5SihzfbUsm7oxZCXe8AjSulItkBkXlvSESG
O85hVCP23d4NaBdQcZ1T29467ojS15m+kdVvgjBxS58tE4yyjH6lRLcklrZbHTAi
15cYLxokQo1lxnJjKGbw/C6IRk75jLzqLEams9e1JyMlILSl6juogJCB6JpI8lgJ
0eTv9MLuFZkD6dGFIndem4B77wvbI5DBbTsvLDlmwTcXyou/GFf2Ezx7rZpenNZk
PM0ZmAZ40RBigMYJWe9/iM0AcJBjVofA64VjsN9G/umJBJjybBduEPYX9i9lTCEZ
VkLyBviCxPMigMjujinJwrCbvSBaBhSJTudB2nJBF/x11kEzfJLJvpmWcxrtKqy1
y5Nca3CRuYa2X6snEesVx9C9FiZL805aaCvcZtdieZG1KSO+ksxy7Gc6jGWsM7s6
rnNELf4gcZ6BuGCGrsvncJbqL4DiPTopENN4OTVyRn0vPehGwIeVDyCPvoyYGxtE
8RfV4RPCtRy4k2ruPTFfhb86Ioq4Sr5/cUL6qdTXgMBYzVX7YoWpQbn2Ov0ACB6o
5X/aTf0HPJKrtMwIn0VohzvHcD31NRhUWStkggTCra3xEmRel8L9lDKysac+y1Hi
1F6jahlLJDJo1SdmoPaNJxQZ75BB9WypFEg782pg81wWVxpdNIrEJLUIjnhd9JUP
J8LPfMAtLZsrQYiYTneiOeCLJv46+OExONx3cfHUMadNzJEFFuuXIBhepkb1Fpj0
OmV2q6p5/Epb33eOXqsLvhVk0EMIUBW8qmj2yYx73rGo2g+Z+PPFgw0HfQ0peM6t
8oScpbb3t7s/m8PwvW9dt4UubQ/HDsmjFHVTW79JBRNp8BzJ/BT9rUt5s6zI9jlY
KcrUVjJwxr6irxufHOVA3NcpYvAupqC82eWMmk1W6BLf7FIbRjf2VKKe1M34QStp
JfFK14H4gV9/2w9/p2Z62uw2hIXjZYNORxUgD8/RbaFQc6h8iI5ZamTM068NHGW/
8nzQQX2gBZ/GJ7tIYLqDC/gO2oHBrgKNX/WkdXBke1jXBklR+vemIPIaYT8X14EN
QVd7l2lDs4xa6JRD724MrxfaHiYLIY+wfmMcTC0Fm0VWlYT3IiLnj2SNAzkNGHuB
Azyw9678kHQpm20l1A7xv8bXFGqp6S6R6957A2EUnDnQEjDS82Gcx1uzATFkPBjC
1W0p/RDM11pBpxhvRI+SOyzCHwqfM42q7/1iMJWE4CaFqSLvWjTkf8li4V9Pxdw5
aizCHm393LSS/UNOH6AL3p+8g39g0liJ60F6XugSUFJPJvuQwpfMTHpyvY8voYsj
akIWGf4pPRx+L3uYFz7+oaz6AU5Tis2htCzhm/s63zzPm67ZbUZImnyLuSBhosN5
g5TAoPN0Bs7KyHSBe8gVFQvveRgk91uVdi1n8dG68tnadD+1DCNGOuUI9h9Saq6h
DHbjmlNPGjntZZ6CtwQXYqhoGNVPP0osjrqf4W3rBZZQEzHhvGLpp0Z7b2SjNqZL
SmSjsm4YPq3dVGGGx+/OjTZfv/JTlqhuVTcvAgWCVEl+GAwhveha+8snzg0yZzOW
yy0qm2fceOKd/ZygKabK2DrnbKYGYg9ekCeRADa3yOhrxvC8d4QxLB6AwmybqzKl
dwoY+nQKQoIFM2jaCI9d6AMNdZeGTSTuKa6ydtmjo4hCzTJe+KdBg30Da7gxsGdP
fOsVfjdUGDXBrAsE1P5YNTB5i1bn1vIu6P1h1gJyEkfxri6fwnmwMkxF0hIhKsZV
wRlBRRzEFGObR6B5An45pbOC/+LoiZ/9UDqrL1tH1AiemyOpqiqZ0D6R74zmzcnE
g+GpxXgIhfE5OhJuy3gwakCK6LLw1QwoXL16sVr2I9MSpeAb9jzvgvRmcWlf0dOG
/ePaUPNXb8ibj492W//XRDIAaH6FjwNWL2A2Mxt906kbZfVcOpl1pDIh94Sfa87O
+RCQ3nP0txLgGvOIZlWmK4QFHEQRZbYtyPl06g1vh4rn7GFieqwZZPzkOW6SOcnQ
pLVjM/lNytO5BpMdVRgUAzZfcbu108Gfq7aKTW39tDc06Mcjj1HWtzV5vs6i9hxG
nsJW1RtRU64JVw90RmZqw7VSrPglr1d4RGm8E6rttrKtVR8fSFxzkExI2vf6JAxW
pYH1tFxF4ZEsfnPhUnglOWnEmPc8gdM0FHzlItVQnOBpNlfSvWtsMqrEMLuZ+1hR
aRErEp73QEkYk9olDW7KhUXCs6ZjE2WcExutzwfzG1jZpNwFkAk6RDXpHgsfbSqM
hBbOC6KYg82cZmXqBqtneqPfSxTX58JZbBAGk7TJ2slnYztH2GZE29goMf8ZpA+3
n6w7lUi1e9Xjg3Ea/IxC763BOWEpxoc+cYcSpUvAxjfqOps/3/yrTICmEE248DgX
lUSUH7pFkEFewmAT9QA7/qVj4scTX3z6DQjpoJ35GMasFDBYjqV3c8Rq/8NNhlgT
l+AVYWMS6COzUEdbSlQz0a/M7NQfM0WbvBAGzcwBBvZXVbLiWboI013q3X7nKA7h
qSPF/whgL0O63I+8FSHqFaYyavnJARAm+t+ATzU7UwqUlkm7f4lrPVehVVRW7eZ7
DFjcbPsJW3aMkb4luc0jXLzsGMFFljRawbqP/oeiwa3Cgiz3OxQVETyMrd4Rfvp5
xbt13tdEF3MxJUGgfbwk3S1jRjP7FpJcIpjO5YuCFJtgTpnnOPDbSE85IJl/e9/D
qLYaeLmyq6Q2DpuAKy5VpEm7T/0gZnlenCrwrbBxV0fe2xw10g1g06Gt8BMV7vW/
LXN3Hol+CASqkgd1Yo4tDqvPhMEK2H1cJ4or3Enz9MLGw+59a2LA1vISKp2RHbfb
GZqe9KdjuIK1sYeR8Cq53JKA+/YRW1qFZLarAV1j8B8Si7piuDxFPpc8/EEfrwEe
N1w1Vak5imi05XZLqrZW6OtEfnFXBBERGESe6sz4CEZcUhG/Cz4yFhXBttCPAr88
akknBh40kzWU/LDysEAVZj/JbBb2zh3v9mrd+gMVFssusN9lbFeg4kgxa91Sba3U
zECH+bIVVAMAbz75lJepSTDpOeNB7JnmJ/dlIMCHuL1u/DOOo3JjWPPq43ZRXHnZ
WiAReu2Q6NbEWyz0rUZ6Iwx3L/zxkE6sVkCmxhRxFpdDZVOPBj6yCGsFXIwB8Bmh
dJCvWz4vWbfyk6pXRyq8dtMLu6dkEOzOpmeUKk+buQ8bbnYumulM8flGLMYY3Z+I
AkI9m1mftAkamZvvtkgq0GRjXRijgXZ3UKksw/NwPt4+Bh647v8w5I6etApjWSQ+
e0GgQlaxfvx1nv3jeRW4iYzY4WWveP4XbgyLnLM50m7lbJprjTWxE8/u7FEjFlTh
yGLlyPUVVk+2aqU5dvGjrIpE3gUqFyM9VLHl2QhJa/JswUhHRl6z+/emIZqsP+/0
fVmqUYZZd9Cu27iP+cISviNzaqi5J+VUareXBcxFlGsy+LkJjv5HhfQ42Akj3q4j
hYn5uLOpGn8tSIju17sqmyMazzy+fnQmmxjuAP2OIe20E00nB9zURV2WG9EHB9vD
qKiCDomlcG4yplm/lx0740mwS5imQlsXgv9KqQRYNyvNpBir4ygvTt20utXHVuBx
igM8wZHm5o+/Ow3mjE6pTRBOUYq5Wdi2lq0A1iajsH7sHp5vvl8AIYq8d/Qrdvrs
gK3g3mA8Tfx12wXfq3NS5EXfNO0d9cIZbm/KZ4tWYMumuv9CRQh1HMKTNwCfehtN
Rq1M4uf6AVGknCGMowRmr3JGFUmpryHgtgxYPinyEMP54xAEAAw0AHpPnPmdJuR0
BdRRD6wfCa7ko/Ulg0issOdz0MrNYG2FdMqPY9FRmNKgb8RiMN8fO8uq1J9NpKCe
yP2Bey9d4Mtg+lBBwWMyNkxdZfj0ExZtzuPAednPz4zw9dbw6sS/Zm1x7RBjNPDH
IkMt/edCiyR7SzDKvsNphKnTkzX4WHZVNXRD0nr/TQM9lefmGH3xFpgGiXjkrg8S
G1l9xeD2B+Z5dT1rOdm/ntygx7ecOTSr1WmJnpUq8B61fDpAcMqql2BMK8W7OzMz
ctXyot6qnJ7VFFVGtTAvSN2DPdw/xVWp4VUISvnW02nkSCz0kn6mmtM1tleRO2wY
mNiyZ7TP/9QNPgsa2aW9C1shDd6JXyzBvQyKx9kdRPDEGi3WVS+AknotZUtVGvbS
n1oKKnDWIqO4zjIwEB+FL0GZRUBniU63FI5dEUViVWsoa3JYll/wucrjhBORIZtX
5pJCVHY7N8BdteGM0+iOAwPp7leS30TUEQiGmm81cvcKTtL6WSVHBfHW8WecPBbj
KfZuQLNUr9FoVHO872QSHl98VbjMRpq54JxgGuPRgvRWccXY9Aw9zmr1AqKo76wC
rM9FVx/TWLr7xFdfjUsXhbj96/0g1JMtw7u5UTac+f+hB3I4jSYCuHWmx7EhgbXr
eFAzkkXUEYrZM97jqvhbtr0csYRmsZmTfiDuQ6Z9Az5rzELGI/VSXGWUncpQ0UHt
Y55upPjRHfWE9TTX4WQns1gIQEEKQhi22Wr5/FV1XQjnl6gOPVWJOIsXmFp24zGC
I2Qi/B4/DecHi0jD5fXer+e+uhAi04NsLfhYT+ip29gYXwJw7FgidnEtOdN73b0n
LyMVU2kQDP+w6/31RYzKuZwWb1hvQf+VuLYhDQ9uAO5Nb7Rc9hTLl4D3N810mjqn
7bcUVOs6eqshEOqZflWOtQMFbB9V0R77VUWDIQ4Gj1KITzs1o5sOPFJF3kH2M4k8
q7StiSBSqUdD9RsB64WqD3W+YEwpRNqnnn84xw1KJSqnxDQNdq+QgOzzDzhc7wRp
n31R+XWavDEXhAVmOp1EVGEfhig5eZc53blKTXolHsjFqmyLFe/MpF4nCxdz4a1t
xmJZ8V5enBnZkAnC+kZhVmQvUN5rDkYZsYUjwwN7QalKNNf4BBXYIXPQRnoNnA6x
MSs4ELtpfNlQbp/ASkrjl+WMWy/6bCfF9fhvOi6fMfcR09P3nndtcMoyD8gvBFAA
8OeNIrg8uuXErNXD7uX8asfJ1ZdgDliuVSmLyiPkMuir9IwtekB5w5qMkowUvICL
7qD9grXZ96thkQ5MXQylGqkJUgQrR8CHKuPIJeGcz3Jxf2nHPq0Baa2HmKnzTvpw
058Ji+awFfHgo6tQA1nfeX7Ow0FiUQOdIzgmlra6/9dvp0XlhDb+ZD/dTrDyPg3d
xaSBWk1+tT7oY1asPXW3dOUIZew6IIutXP4gC0WvTzNaWSUJr4MGK40DtBEpq9es
gPO07acx/kUqu58eTbLcot4rOpMmrCbRpTb6RQE/IMuMJ6JpBvpkD5dfWPiRiZRJ
zQ7p+PwDCsPm3BIINZFlnhWu7xzFXc2tbytfAnYwRtE1Q0y1bd6KcUid2VXlXHSY
VxkQvfNveFw1kwcTTGdHcz15smI/xZk1+vbHYrOAEOZTbWzkNtn0PaV8N6PqrJWx
vuB0K2kOorb1irlJnMws6GT6GFApaFEpBdvMvJuhFrZqicsqVFMnSW04nrylk9sn
5n80CGhf2SZXBByuhP+0v7qS/5xud7IK89gxrW/4hLCDnZFCEe9KcP8dPWFzkvr3
U4alsoXNrCJN2Huvf5HmYGpGAs6w0R8AiH7bV4pl/zwujKTtwlfElfLV6R51Mgk+
Z4jkayFFaM49lj3GH4E72RO+Fn4TK7hSLZQDJMSTN35BLERRKkBOPBbA2MkCDfJL
Wz+8AuEXf6kXMt4CEfdmVNBkDj+QpMecqyHDUgRQyMJWm15jBE5o8ob0vvQ8NQvF
2ZiCrKOR+G8AytlLk2eRW2Dos5kORtHiJ1BJBv2+5GM3/pqDFyVBbVQGro1xezK8
Fe+uvfp0IsolqYHzyg7lk2UW4ehnnnDDxmIgER9IN8IWssMoenYxkp3g4lsrPUgM
zISOTaaDtp5n/PPvqHkNtLYb+Ja0FpmyuYxiurXEtlk6xoWl937ITAyv7bUwEhwg
6fQUUQOaT0CJ4+To7XyOkhvXUY5bWfXODGkyX9eZ/GNjrURftPzXSOz3nnue1a+X
4PcmMCrv4a/+lN93HS7o7tdxdpHU+iugbsg8TzpG386HCOmLB9doRdkJcIS6tY/A
mzh1vQNGPFgYzJ+0DCwgbNngnPJK5DSfXcPmcGsQVSACU68+ozl8pj0YJuZDtsGM
WhCfWxyt31y/l32nWRAG5cILX3NUFVQcKWTnnSKI7J2fHqO6curJZfmHXj1ljoIq
jHL+LV8AP9nn2xMkb84zV4n+aBRg67RHJTftuvsWFfkmdjsYSS82KhA41/06n2MB
LgQZfUevXaNnsgqPwcOFR+pALY4FWEYE8fH70hO+zwv/QjD3aa8hyLRAbY5FfNGg
ogIe3rDutDmUYbsY/onmbCaOIPE57VfIEBwaExHdYdpXwzyFWDSnyz08ILu7Slob
lwkm98pbwS5bHDMQywhiGoG8TxTMDTOFVbrcPI08onSVvIEYOsEhQMo4HBNWk2Vf
79JZdsO3MKqqh38bVaYpflWR7uZsKNp7VMPwfQebzaanVfVVnFMeOpH4bBeAOole
5FHp2okbGMV2CUEpQJPMwu4WFCYB8xqviQNhAipaqM4o2XOLJrvwUTKq+CD+sr0k
eABVgTn6MbpcOH5u3n9mcJTBchgdg1CpfCpgkImY9BXZoTRx4k0S6ioEEcsyVKSt
0SOm+pPshwBTz55Z2ZJCX1NXK/g5uIfROnS23WKcDR4wA0NIMMWhi7yrc546EyGT
2Gg2hMjj/k+FtCmyuYT1u3dmoODkykG/aQyAXf4T4M89Tfga8SBSf7zgcJDFI6Ua
SfSrOHjT4z87Giggh3PBCRZAYizfRh6NnlLcZrTtEuIbFlFOiGqbTOT/YNjzeUyW
BM08eSZEgXJQLZu39g5EbWgrwerAfJoayzjFFJUh47bPWWYzawuODaIECUABtzjD
Dq1eDrJXq4/rquubpof/Pqn1aWI5mKUx/LJOMVNCvyCdfVEEOse0pEnVkhDOn1bp
v7HbV4mFc3x89n2vEu++poHWYGIAkKS4lxaHbx3W10b5ijza/4nboovHtgUhA1Xa
mb1FuE3XM0jdNFvx+umGZBRgTKJ0RdXGi0fvYhl3cyFo+4K9dOXIjuo21oLHnTsy
wZAlAQ/J8F1jV4vlGzw27LzDI5/abWj+Elqj+mff6igqaGC85V4YslGCtUqmK+Ow
hqn4JAlyVKNC5CCs5+XTq9ZpJMhdwVYbb37AlSoc0kSzeNXc8jqCTRnoRnNDNdGo
XS7OtISItnoP1l+IBdgXd0LGfFV7BkQkKa0Pblvik1N6oST6tUvMsCH+esqJRkSB
N617+YzhDFKJX0XNmEQef+uMMjm7UsNBMWcRoAVGuVebA2Sttw6/fYaYy8Ksg7hB
IHJaVbnAvYcCmxDo00XbLckVpaZMDpewP2Dk8hS0QfSvLX/oswegjXLG3iQhU2mu
LN79hN/7RwFIZMbw5oTQFjDkHJyDHZaYr2WreUfnfEglveDTLQdS2E0LoTvx+JTo
6reoO+cbuZr3M/V8SIhSzDayvpIl6c53JeeA+mW9RTDM+1UFY32LPMqyFULhz+4H
z47tth1vlPlayHWTDijNrGWcoT4R1Fov/5sUKzvhTgo56RAZRQ1PZK3LzJ4H4cvq
ryot7jX5x7yU98MgtnEboxdqd5W4p6PgputBgNx+FayeAXv9Siv8bH7gr8RQSsy5
AFVdB3yPnnq5Qs23ndIWZPkDAeCWk/mdKTHRzfWCjDbp77ul1BvMGismv/9iNnB7
JFYcICmNnubkrr5RRv0FwDqBVL8VTxZvItjga+UgkIpfia1BcVu6sow+yev1NnzE
3vwODSIblcgr1yDxFT3w8oajFHi0YzUg/y9BS7BztpiNsV1CoF/WIox4DdoZU0P8
v5J8mZFle21YmDCOSJF7rJ5d2YkyuKsgeyqu+slSLsAnHEpiOqAiL9vZj2b1WZfF
vvhSlgmf4hj55rTn7GqeNUtK9eSFnl+xRMhKDitqX/vLUjD8q6P4X6fPYSYelLsL
BfuGTE9ib4SgaIunWg1S04yG4Ol1zJqEPpl0fRKOh59wNUQg7NwhjwYIpdT0L9Bo
UlIyM5ePQ5oX56r1YktY4FtHwt5cwG/3P5geOM+n4iVx7wdg7HVGLc90YF2IxG2K
9lWaGDgr5/WbsT1cX3drNY+PtpjhgoIna1minaYVUunFzta5PTDgAMofbFoTt2rh
RB3GIFrqmh2IMd7yBNDbaaZrI9G7TVj/Qft0yk2Nr7gFxnhds/B2HZY3cfuPwQtb
Pl8lDxyHgcw0xmUQMiNA/UkGP4tuUIwD+iOVR7Ul7sXWkzpb/0wgFxyThf4DaES6
XiEaljisOcBWEr/+0kkxUiNzXIb1LrJObr2rP6urktJExAL3nWDSx6u/hi9DRW9c
FR87aHqkOGWBw1szG4TOFgxSwNNUlS0NEPnLS28pejsJzU45MblWW7DgNHIpW/9m
ryj0gp0/l8cDetMczq93jpGL1rPWjd5oN4NB1GTZCrtXik2G4u38V1qsuCHA8dUV
Zyu0Eb1RVphmenNpGQ/CmyPGErDnk9OmNHL4sK9+NHMW17AXG+O8ScNT9+eTRSzY
zoCmIoVKQ2GzY8diqYILFhNKifQlBg72u5MGIdmfq3jE9EMqnW/vTnRj9UXQ28K9
mkG2K31jgnc/BqrIad6nnwauECBwkktbKg/Gwe7zXv2aeeWTjk/xpfaaq4M/pAV1
0Vc1haJZC7CaDHiK7TwQlg7JRC5ub/fK+w1Ovn5a9oJVsapK/L3xUrn//rPnrIIk
lle9NyJ0Bep9qj7k/4SjwQoFTbN4CMYPoZ5zo5ssiAVkWbW3k4+35x1XhUnFOIcT
m3XnGkqCCa79MKJoFEeNZGckLEB7WpdoDEjsM5pvDpJ7GSixncEFbFgUUsfTVjnX
p9QexoCo/f0qGIYejKUdTU+43P8WbIlf0t+F4htic1tcETiyUF8P0R0w9DBTmHRL
/Rfuc/ESc5WAMH4MAbPUZTD+2KFhR4XK3TmQwqdd4wxPHt7i8YyxrJXkB1PA6PFE
jDT+Uh7Ojoyyhl6f8xbE1nmWQ4F7IOBtVuY9xSui1s3doWRci/ZHtxDixKOswNRc
eLpLoWSrpkcfW7IR9HGGk8JHkaLeGVCPoFuGu3enyS6Wlrhz2Tq3w7IznzkuENEK
AkvyjfQ5r3HAUahvX6o8DriIOr4ehGbUCP2uHaUmGqMpRdMaZfekZj0+hqOiBWg8
BEcKs9Pjpb0LwanNqmvjeUdI64kq+qZ4CjanjtrCds39c91+Zxid+/apEEtH5vhx
8cDT4Z9qYiSXRvui9d8VBqvdkrtqj5E3qJGKEhvMtrTAwDVMvqWRPY35z6Tb00dv
1BX+vK1/Q4PdfDgKeEruoSYVCJLnbUdB+1j2dwKLkHA4e1lZ2B3hC+iyW6wfr82j
j+Kqa+fRX8rMl8jK2XY70BmsEyyUPDMy1n/Ox1rjPF7orBi12QLZGsuF6daiLIK8
ZZOE/pPxaJiugmEiue6r3jEwgi75FMKB3b+HKCGAvjXGEqNhE/+kCVsWfH80KnZz
W9wY9MBU6EII9ddmcyyfIxyBtQmg1ytxGQ2rKMFBP6rScT0a9/rIuT09wVbX2kA3
KJY15eoP/pEPytVCu7Auk0V+JODkgASL04Yxe8kPxtsJ2vevt+FIf8mTFPOI74tX
aVg+Yani2aUJ+DaYYfN2Fe3SQA2uDRKRj/jIioz7IGq4lyo1fb2NiIMw4nihtHOT
8FKAkk3wcwUdiFdWvglDLmmorWXn7hNH2Y0644N/bdwH9TfLlAQuY+MSZ/oZr5Oa
U/ILsZEGlu2xlUSoh536HJS1QeLGYq1CKVy0pPba/YiDy3VuFLsZMDL+HIoxrbkg
MxWBWReyP8HD9F6j2CqC4ik8NqpN9SRgkY2WQBbd7DILkCgHP9jwuPZc2XTZWqoF
FwWpq4ioz+WqR95BjTcm+wdDV6M383bIkIIyJRMRvRu8y75SwQclWI+eJ6Sg+IID
BkYz8VXZSlbkgQfH67XUq5HLegYSKOjLuFS9FNpexxOEBctsgHS8vP40d+kYuG5u
Ia6nFM8jVaQoXjAxifoYEv5ZroivCFQERBkrwIWFfWYOkrE2sXlambnisJTzXZJq
XNAu1J5B5a2emu3Pri4ozX1vx+ewYdL2rCEbP3yyc3ScRxdd9Hr/MBnbu7ffv2yN
YfmjZj0meTbA8YHrsdHjDLnE55zEDe+VBXNZJBpNwJjT6GI5L5We0XOh95KjeNhC
TZE+BkuXmZmFpYpLrItN4NJkfrRu23kacofZGdza0JaUavtIfiGSn2scaGwUnftx
jWynWA8ofvBMv1dUr9byJrEDwlu4pg7G4LkfHVB5AWUAdiMQ/BescF8X7ULU69dJ
P1AOXCEXxxcUUBHXe6tmUA2l3Hd8yr9y6uub9ZQ4KCvtRG8uVq4jM8i/YsKPxv+S
LI6BLPNvMOAmTAJ0TFE2cLc7p3ZSp8rCPUEN/b1NqG4ivqeYTae7y0aCyuPgwXrL
goom047W0fvkRHERohxMIjJXgCPYA9P9+y30Fq6/9GxyKs9ZlGgKGqviJU/EEzpS
wAOsOoo9rhnQx02nXFU+23uWH/sw4+hrU9/kKI0LjVkW99j+4rTIpYLvhomD9LVD
QSBX6H5Z6lynbr1xMk4na/Lxgng24ANrCa/WsNTvsQeiHQKMnxhvwRTgwRYJaTEN
sOqXAxC9MdqiMKaFpCyDVOq24xpET8y1rOU0iHrKr0y8f41Y3ifP6+wNR7MjWGYX
SpG53MTZy4ztpm4ONFaMYDYpbHqUfbw7JCnI7JVZzNV5ySSgqroq/P8xr9LAOXJO
869LQr0j7N4JVP4oZT6K00Cdsw8nmxjp47fUa0qo6CZ3JCGWYTBWyA7z8WKci6RU
5612vk/Axuz1X3D6b1S535Qj0wVu0YstFBQfKXDGVtvf73t4OwMwMH5ZOMTYbPYR
U9Nax/VwmM02iLRTvHFPZeRZcmKDoPjou7wumB7Fiw9yDScmHm7kODNLDXmnGZ2c
w+HYlwsN5b10P9nu82hX0LWmCKeOROIZD7b7UqxHJUwq6Qa6JXtwV7Mz35eo24ge
7GL2ZdSA4Nj2SjotUNkjO9VzY+CqVsLoGNqzobcW7+eSmMJkslXrlBewOAZVQr/j
UGZkHILLa0M896xTOo5zb/VYK1d/ke6AzOtPTh+CYlft3QZBftTtV0uFTW8s5YdT
d7v3bMr6xm1tnJci7fpOvjEhiV9Wj/gHxyHmAJ6ilHx+dEf9GABLUXaJMfPucyAW
GTkkaMKFDFbs/iYyBQt/JjuzHAuYmB8sxsqmqDC2UIg7Vvsy9JH/r+gOBTyR+wk+
K6TLevfAJ83k1Il5lLeXNqO+nmldzzpYeSAsI+KuwUKil4qIMGmjRC9KYXRfRUNz
ka9g0Hfc75AuJq+R7ui+vPVtnPn5GjMPzsOBNnc6CWLmle5nGKYHzz0tMQSISoIM
F8UZrlsiFM9OKd1rXmvXX9wrn47SQNS0VpZGP/3bkiGWsMMI48IRl2q+NBfuP+dZ
hHzC5d5xbd6aQ8oD6TzwHsR3PsUV0xVaP5Dk0H20cWGCxrfgvlY9r/Lmu5r75he3
QudybcZthfQzA0FWXj4QqD7n1bIo14PKch2br9+KrMWTpznF1wC0mYMmiyk9fuvb
N9Z1vKMbkqAjEuPK0y+ewQ5QrS5dkTLB1iaS4MqXUH6YmxfPANX3aYVte3i/jSWW
akK0AappglFIKVESixktPdworCbTtYkRg5yyEpOlBYCvIX1jqqA4FG6di9OPufBQ
hlCOLRKf21OBccZCFlz0tPR20pweE8T7raoErJeMMeaJLjAu+mwjz1+nlu5q+Owp
0C5jQnxUJzlfrhph0LUqoFys8D/iBzO0DjlFFYQeIE9pShcaVqi5DtHtj/58WTna
PEB0aMM3be4eXkFKVM38b+kyjtyRdR0JwX+wAzMdLuerxVWA8JqiqDEQuj1Mvep0
dpkZ7ZXD1NWPPT+3B1UQzwr9Ajy+32j2y63aLvBx7fPRmPgsHdmXjSQoL/7TZv6W
cNGUPRTHvf1RnRRCaQQ/hZ5ThyEYxsaO+W6yZ3cFExvmTurni/NmU7/jNalp68jU
0CI03FW0zltX3zRMixHuNc/wB9NsllgQDXXiUg07IPWjuvcnG5onTPCpwyO1M3S1
LYU88Ly3TkZCrZfZIdjsQswWQK3Jazt883bECb9EdYL3Hgz0SA/vhADiIFu8EIPj
qXI9O0qIErR5Il8uQFQNnPkOEro5PzCtD/pXZCIuKy0FeFlc0YyCHTgoWr2vWcP6
9Lw/7Fpzivi6KGW2CeliUvfpQa7JfZfb+uVRCBI6Zn5vglvcJDoXOOYnRF6U/zBO
r9FVaURgyehsjbgcU6SB1E3HPIEulerzqtct8pKZs0X1Q63GW9LczSzCYp/UytWq
+t9LWyR9m4XLic6A269MVLaKxjsqQPszxuA3j+jHeCOUmr/nx7bD2pkqiCXfnNnj
ux/1rjsFYABxICcpTJG61D+iCNLscHObVgPjhM0bypWg2+v79i5tYXqzeWXkAUYZ
SodsHh88zbN3AFD5n/7g2FSrpGXhf4mbrZNF4DhNXxHZnDzRxKumY9K1vGMJd6kS
mV76rfGV5YjCXm0nsZq0+KfbLCsJHCNmiwepREkiChVhljQd/NvUcQzKBhjU+WIt
RNXOmDtBTGQ+lS2lbhJq2LIQAJJQ295ksEnevFVo8uSBAlK05CLwOR0x60hotCPQ
tVsOSTFWIJwgZbTKnG04s9aAUNmwHQf+zW0EVFeCbTuvS2df2u86Sgv7iM3QBrWF
45/IK9Xz98mW4U9ov/tZ3fbs9udjoT2Hx9ZlY2T0p95VPVxj4sqCPfOUghwrkxM0
KNzBtypBC9pbvWjA6YXDMp079x0Eyz8+d4+pF2JAnAYjX2gasSUawyKj2yjysjrP
VQNvk8glsqI9PtB0sygeYMP8hEV9uuM+Kx2oj5vGTfaehxEtiXIlTm0uCmDVwMRd
EvnaYvtJvK1l+Kz5TEhGh3TKn4L0KosSkk1GdvxcjTcFUAh7wbOt/Rkq0L0Gfee/
LmZ7QtjPm6uTRf/IrQcnoMgbIf8LgBscWkcQy7ic4hA0KG0SWtQsldc1ANn+zotp
WNdFpQ3RJQAz5j73AHi9P4VVEADbPD9933ZLT5Ql5etQozRmwa8XPDQjC2/H4C1a
811HTIwcQszv7umSWdVlNHz+yGPoywqAOMXtsux+8K47GOhLTymPAkXl8Hd3J64F
1wq23ZzWUgBtUaZrQtvtRRiXKYTlR2MwkFS5VQr/m0kiv0lVFkQU1C4LsODjTGV0
/Jc5vwHaIUzddCnHWW5l2Iq3bBXid1dl3dZw4rJaC3IV1dPXuLHF4VLIEspt3RSS
oKwVHJKfPkT4IuXIYs+v7E1IIEDlvJidNz2ZOVKPACiJ3hjMwMJathJ56G1vXpBc
oy0qo1dm4DOjTHhofPoHuNzxaYmYRQwB21k8e2x13+CDI59CV9Lp8zXIlckns9kC
r5vSYWsLnnBXUxZu9xG1BrwrAMsxl4sZ2PhlkB5n3aHaYxdo0aNaGhDqI9SHwlj7
nEJm1qWzQceluEA98SVcZ1A0TuCD+5uNKJAsaYQyrtkNE/fT3HV/ZP/Ck3xut2MM
oujAsy0psei1t+5keHXMP72j4i5bHrY6EVJ9nCCuUZ80OJ55uH7koW8BlYYxnG9o
uHAlvDC3gZESaL7fS19mrD4Rbq55RSWd0I9+TexswK9TcRWcywOJKAQKfDYFA+y7
CDcMFRCHgCIBr8z/F1TbYdEqh3lqySyVb2l/KaKh4vPu6pmQIOSaklLi3XR91bLS
BPMe/CLM+I6c+T83ZRrV7xZd8FCdybMS9Jczbu6pRWTSK6gGdLGiDvc8QMosMPE8
JJ+sle8XPMDWgzOC8jYLd6AyKUjpJpNxu9Hah4tr++Cg/KZVYJx+KPjgBnHuHqB2
7+OeYHnsJAr93vo2BN/84P8SHUqFlCWOHPvuIj2c8RHmjuPOq3kubXO3+TugF3kD
vMlrB2rWyyxCg4UN54DVR3XqaVcvI11KtNx/WZNeFZDWaTNPzB7sCPbSRwLjEY6p
Ilm0T5ALGIry4K0OlqM2WvrdZrhI3NAhbh2TxuP+eNWu1nQ/McCFypfZCAHkfACl
s8zWfv5W/GU3A8X4nYcnwSSh+aAxi0SoCBPunU8soUkbQpXLDvOEwJ5negLFcDwn
AJEVi+7ztfEBrXsJ0I7cep4omcYxnMXvwAbXxqt+ZBlcQsarumZg2X0DWaJlmMlr
cefeyyRcNwzLO6ON6yf4qtXwvPl8EoFzyKZ2MVpRxTKrUwA4DvvCtOUJUsOEvIsb
SsDmvbmZG5lAHhSxstLJY1N/Gq0giORx3QHpD8HtbsCoDwemV27VBPLdbyUz5SYV
Dex5vG/cyiWqIlVHaRy0kktztmqmam4+BW8JOwlS+LpQW78jzKdRheF42l6ZZjfg
0/bkllQ/9is0ptqnwXa4Z+WJTHRALqmgHmEn1LYpDr2DEX+8nTpTLrBEGN0O1nDi
aqyEWL77CGH9YPy0U91BIbHzayVkcUJWmV4FVJfwFKTZCXKuzbMGqrwgRgewqdJf
TXQRDuuyv/YqzezDWVFW7L7IinlsstjY3GUjv1Ca/mi3z21WkThuC0zidTrT4jY7
GjyhMOK8oU6+c5e6UBdVrzRHkDvwjpMCw9U2ZuwbsMVoZH5pU/5Pvk1VAmscjErK
Ol5UgER1M5CU+l2IeZV/Zy+DrR/BvSMJJSK2RS4j4vAdlPR7VesA4UXb5ACSh0ye
BZ+XWUEbzevDddVPZfKbLCVxw69k2QXGTplnIxT9/T7SyBIrgKICCwZJZA/7LZGZ
jZ5EmQc8O6zxxPCyOumpL3dR8qWcgMEkobEshY+MPkAwT6sm6pfvXecf5MXwrjAn
oU0nFUCpL87Wnoxa1t9KY0s0mzF6YkWkRvMEcSLQ70kd67o/TpGiDJB2KM07XwWx
foWE7FrEGz6IyPqQqg13xmLlMhTYGbbeNc0X+nntxqnrIYNRIUiMTXVU3F7zYTpN
cwUumX/6tZmM9mZ+0A5Q3L9EDrdOa5qdTLbVBt/Nv2/e6dvhjZSpZi7Gw1YGdGvl
hjMtnbrKSZHF16NYywcFOF6+lfFlmIR69n+PetC7MINzN/s0HWv5sKzDQZ6JLtCV
7B1JLwBbklpFVciQvbN+1I7f6/tmhXfzbvRDqsb5xQgy4Z63MSHLZ37TMQDOwXuj
kOjPA58lQ22vUrfx7q6VwOYRqv34KWe0l+D07FTwMltHLs6Ps86qblnmyv1SyOf+
qhiGGNOc+eGcpkmLLCb6V2VnRtZAoWleYJFP73UlbJ56f6adTbnxRnhvxV1gtZOJ
Bg+woZDOHxf/FdxhZFNezRGXPtuWsk1dTFuLksL2Z0iOdWjZuwxvhooXlWu/K+jf
sNC0Vlk0ld2DcRF1ButncoNgT+2muWiLi/UaNitgjOa7iDfiQt8KfxhzpeWgXO+0
e3JaPwN1t5kFvttXvwzKgDUE6fbcfyhM0I9lmvWDLK7S0IUVNLIn4X2449YTWwt6
EfsSlQeKb6BUd7MTh9q+VSewDSRN0K7LuvAAklC0E1t0dVgAUVOH5sfKspM9SfKj
EMtF8EUAFP0aHYEjZs6RJL9sBW9FUBhmxkbKegrQWDoKIjTBF2c0ryiDQOfgNEFq
Zx571VCFoooos6cIJQyjpqhDbd5AVA4y5FSERZ8qyv6VBbUGnkufAFGGwd4OjH0Q
ll9Km01gjRVFhdraZp93K7GtVYymMpXB7DEkBCMCVbSoEZCR1zcPJiIga/fZoAG4
7r1KivVh5x/AYV5w51GkpoS0jNTGi/G5pFXj9y932DaLMplTWNlXp1ssTmvHhof2
9vHzcvaLSjkCiwclSShTW8p4DhTHPWjtTzBdaampPjxOWp1GmwTqa/hc+sZ/Dkvf
nAOLl7/7tR6g7+YYIQya/RVYf6K9rswp7QzAmiWMCAJS9UbCA5e+Gm53cGMkwVww
t0csqhDUuw4JnuNFMl6BnCW+8nb/ArQ9jY2dYSBNJduM3fUCe+EL9HpexsjdmXD/
3eqDlOU7sEDCliomMYid/hBvf4FbNaxzEKTd+OT77L4mm/I+k5fsrBYLPsVU3WIE
/hM9dUka1Fs732JmjL64plMA1s3PFtY6DEkAXdT2ion8ZkDp5fdkRUrsFQqsdkiS
Zibd2FPwBZ5/BoOQWIr51ffg5lEQ308KBRNusMcdLLr3yjiN3U/9OCSsI0kU0KPs
3ZR7RnLgcT+UXwO8Ow7rAcKBNcvWFhr5vQVW8u4ftshmaSCMs+6drZgOz1qFwONw
xupjwVbJY8eM4/JeXFQ1TwPA5y3gxuns3YWZR5o3+CRBdqqHp1UnkSBK3Fn4sqKb
M7bXitfcRNSrWCDtLGBbixbIWiDywGRIIW0xAbK1mXwLQj7kYY0lPkXUF8hqhybn
lCO1vlPBoS79Sm9Ea2evSw5TQqjmviVM1JdOXZ/chz9pyqVHkIPBUr+rjBV6t+s1
Hl9BHqNlTXAOB0uwC2mJGwUR74+n7ES9QLSi1UgxxD6pMWQHO6ncC3qTRRUDJoHc
1EiJ0X3pnyom0A1ev9uw459FP9K4kr61+p0xo0rc9aF0u7ekv3XeiNls7bLITf8t
25PwSkJslMdT7dCEhL1qsj8wWaX+YjCJ0d4GflX6MmdNFBBqtXENA7bZ3WetKo0X
tY0VQAU1eLv859jut5U63aa92au5OEvkGVAWrQH7EMDn98qbWVSOKNVpFHFdvtq5
T4HREkO730VcfG1zppfeWsPLXCN8GDlfdFBqKw3UfXqPf7owAOyaz8Xn8a8/jl9I
GOBKtrw2uQyI7kjXLaBi8akrUycvIIZu9ImxUad1dq8JGZw2E5o5yFJUT3Q7UyTg
VsWiHoD09xSdGhx6b8DV8+FWINXw7cRCmaCrOVgS3lwiPYPw/bmQhzOoJnrPMo9K
C4Oe0HRVU417hiVHqBCabJ1kphkjOny0ROJM3W341aN6NyHfpNQe0d1wBHXEgqFs
1ZF4g4kxkZxqxRFnwmuGuzbFGtmidMaeDyZkv645ctL4kFazJB90Zdh0ddoMH4l9
9eaLpGOaVZqPyMXHZxD+SKiZEfox6RXbJUR3Nen/uEJnQIGYVYXXHXXNcfwW30pM
DaIpsOxcf4x/m762gvyhLhHpey7e1LDAiqDgAIwHZk196ozANmr2TCSL1YIyQYWj
Sge13wj6niA8dlSwYDs9Czk4e2vVqrshrCXVnmGyphJGLI7WnlIkDRXBxbD1l7qd
qDehmCuERQdqpGACjX6JFITF3pRItKeVl4OumtjiTVOVUAm4mo+CBGy1HU/cBnFM
MrieK0nta4RqyJvpIVdtEwIYELJB8FHDDRktS3Cu13pnMfEy8mZoMgRKjsmeVx63
33ywr2Z7Tk0pNXMukQYBbTrareq1RL6z8ysc/7+ATnY8fpxbMOz96SZWq2MiGkDJ
rF/KULLq67tFaGvqCN5MvOkfBmGU8vZuUzsIEaoDjypMDAwGZjgkLXD286KzmXTX
x1DrhskE0tUuP2ta2q3v6kcw3BmBs416Up3KdlEZR3vvG/RdIIXmI1E4SFyP6cGc
U660hWopPLd9SWYDe80OlHStqJ7A0GtZB60ZVP7QdfpRZ2324x2rQyIHSCaffJnk
T51R1D16Y2C5ELMgxl30AhREMk5iHgqy+Pls1BN3HkaqfYQjbhKL70xcU/fiXh5P
HDL/H5iUfYBKjUpL871YcaCRF/sIbwY4ABwx0OuuupF3oWvOURFsthvEMzDWNbiw
Wd1nwpNC/oSA455dnePbP3Vy/I6A4gDAnfynl6hLMAbRvPdx1iCdbiZ2S2xnAR4Y
a4ubQb5gW6r8JLVHF3ilpph2bNCtX+NylJhrBB9xOPiQR1q3wc6Sdh47itkp0cv3
wOIZHSRCvFnht1Wu0JsT3wbPojvteYDbnwvyveVn/cyUSVLg7hoMXnXKNa4YKzCL
lEkMUEpNxmHZQCuAaVq4kwhk5Ys/X/+x8UysAgnTTioWCdECR3FalyvWEauBwo99
+DdEHnT9trdeD+4hrc0/7hEktJDvPomM/Nq6mnny38NgWmoTVEJny5otl39CWwBj
2kV6gM+DrRTD3V+AAufmljGLGeZJhPHzLGVXd7DRKasBjn3UFgX6SgHJijrU7Ekw
baS1umkiScmE/izx5QPHiHVroeYaWufQa9iSELdV2j8uufmmItOEZv95FGcaPGvV
IbJppG0dsVhnXL/kn3Q1yJ/2/3HN4Zp9ZLTRBCpFUQPIzKHcUdIdcDXahjkyGDnJ
NqI+YVdYijySUvJRnogqx5eJi7cYFO7+sRp2T1k7ANWbh/s6R8pxNyj8xTYW7njQ
XDwf7PywwNY/8CNQfX6iMVXpxvM6ViQ67FCaLJa+QKJ2BrwXyacBBUVGHHiWpP73
YF+YIJ7sL4IaZME/YaVspOvxpe2SkzsAulNlPbcJeZhJnEBVB+VceJGvNWeqZaC6
t5JI+pJxqvg0Axqy8CrVvd23yat2btTGovT7oyMX4lFL9m1x7MOEzRH06nL553Yf
Tiovbxk+K781zHkinCU+zgLz1V8J4KXVhE521tVlvtulP88BH3r3WczaoY4aUJeQ
cLwJUNK0oYL/Sc8wRxxY6hA90dtC2FMzWubUpei9nMrDK73r2gBN5xRdx87PIkvk
Xi0qSxf8P/RYCKxFN55CvSzxGZU5wJWcrvx/aszCQK5wUonCbPH6wcEvIzcP/1uT
GZaII8XThDcYjz2Wr8nLL9vfkq2pJbZuenF714PQME5pMuM4Yp1UH+R5WW/a33aM
Vn454bhkbei4OHTDmBmt7wP5riKGt+y0KClrs8BjT2Fjpsd6Y4Bwfsfk/TY4zLJn
SLuVcvpu/Ev68WywgyPJKPlddzyRj6mQcL7+TTHwoSi/Jo0wpkc/HpPfBFgPbeOi
GZR8y9nwxysmgOC1MTSActkGERj8zxr7YmyUpFQrggQa14mLLYD09RpKQuAq7H0R
RI0vLOqc3JEMFmRqaGkKUwH9GwpsYGVoulLy5N9/MdT2OO1rR+qoDqK9Kwf79XDe
ZaldIYXnO0nQXgCSLe8XrDYnlKkqfkrjdS+r1cMWEIl0c3UhEi8w+RbWqVL/s332
fxXsAOAuDhZTaxWbPFxnoHLG7Ee6vzQvcYF98fWjHxM6PJUr72hnWL8R7w3kHbHk
kPGzA7c2yRL7t6q/XXJLsCL6LmW+6TogafP4L4XxuZHVS0gQZt3GOvM5EMtgDUdk
K6lb+X8U/IFywYKB2b7p1vc7RQNbVwjRjXreNMbECtnz8EvYZmiPJDM8i8KyVi0b
fQ5Lm00qmYZFgkGzuQQ9/1BfWTEZXPHVJRF+jcQALJnme81BsUf3SnADZaX6q0a7
MCoSG3AGNQ04CwnA2MY5AxajN5X+mu5M1AgAyAQUIM7LZ1YTBq/qK1qMJy+A8SzM
1P9h96Ac1bjxTfFCWy/+UDYLCzldsipPJD4hTSr7hOZPhHgmzSnx3VMciCp/ANqE
kW5mavWWkSFk9D/HWGNtcjjuTmsf47nxBN4zAipAbiEk5KqNGXfUnS7ERFHUsopn
LsXkkBokF5ORqdSxwUYKtT42BhQMj4ANQcEsGhIKLbuaa6VVotG9wge3Ez+Z8OPX
j06SMv0uOk15gQGekXfJ6IUdM8skVtY4vwxceVdZIKLDqom445lvwy9lvqCt1qRJ
P4KwbanTiTWMHweNPwGMlzX30oSD1ALkGu0QgHTHGYKVjKFv95g6F5UAAfWdb4Eb
xJebBRjawAQ5nzurF6M1iY/2OLldu5CmZFCZiY/U9VzKdXQMQ2KryHdHjBelKFw0
I2GjAlQ+Idr42sG1gp8Lczm+p5RoNqfVI6/ZyBAQDBpkutp5TuUhKKuLGn27qxao
7SH9W6Rvpy1xcPJEkEFTGm2eM9AI6uoWkwET0/InsVPdBEj+Ia9t16gXRqaGslaA
4R6idbLsbQ/PqnmAY3dSAo9uTjJISTw0PbEMzqI6RhhtNR1DXTKL+ispjnM3CoHJ
CPltL/khHBeBSiIFPQJTG+rT5245RqfQLDg4o9GSxwRNgpwxY466+uZnWmIllcks
sfVujkrn4AxlejkdQyJuZswLpA5WEclTto6bCR++sVbjkp8mwcke/KqWOZtHCgw4
SgZ7XGYJsm2Jg6Ue5jGHyaX7+vypv7HQk4lA3bgD4a2LizA4N1g0zGYt9/IRaTJ6
KCYzK2SjQrYRF/578+UiFjRokpmphVQIRgbsA1dnj8BuwfvJ8F2ONtxOoao5gtdv
D+C/zLyWBrHHBI8JRItyXv8rk/UQxsdD1tlI8QpgT8MgfJr9l1a/yWaB0hfn7O3a
buMIeQfpK3Uxv6VSdcVe9JeMGeGNsQ6QaXfw3ABnCw/w4bl77rFqCmdx7/MIi04q
508+HEvmMb5MgIFyafZMrwOF+7KSuHJwwgL9vgkcZWGIRXAImdqB2ldgn0dnL8o+
twcxKE+1dk+yiD3cpmbM8W1aGxyXakZ7h8scaTHJBHj+G6BJDKPlprbSglax1Kq1
t6QHfE43cjlJJERgnQJyhX5iTMMxSmxpWNKF+j5fDY3U73vOsmz62pIB67AHxic8
S2gEKK+eGQyJwgVUcn4Fcjb97mTLyTavYiEHFA8+Ee9UBuxpfO4vA3oTbLm0O47C
HwsowO9JyA1DSRgYY/hV8fqcWg6mg9sDta4HuydZkUSTeAxkCfSI5yMmZSRjZxBS
XPDLMLhq051SrCsBiCiwxYyPm/yHlnKvWcjOTyqHeLKkHx2I7ggrGwTZMyXhQSFL
bbv6Uthp7eEuHlbfS4CAnlT5JE3VynUl1LtUrXdMSTFMWzpxpwQ6lKBKCflSa8dq
7qXC4ihrYZuIGP7CMLU4GnosCDNW0tnT+RNYp9pqpKOLu/uiaW1D2/ZDWFwnLMoD
FIN6Aq7/0937wSmjkTVaR5mJhgGP9//sY+QIdOs1xBavTrt/7PGvZl9ee36Aw6Io
KB0N43Gr9xa+LM5POzZZ+la04/kGAarDSggd2CP+JlZW5BnvDSIP0TN/32hDLgvN
ycXjvhtQFzSQGbVfeqEy+GgqMvGdLF7rP1Ljq62iBz9KtlbAjsWoYnCLuLaWjjO7
npmNvzqSod7oKIyRsFVDVY65iHNy8L1J/rhRwd5Qz+gc61//gPz2tb084noJmDEm
2N/Ro5rzJl01HaVWKcx1xukRFuxU7URjFjGGttEM03NpaHRv3mDUY9dlvjRdGNLn
71e04vTw7sjTNCUdoAHy1hirqPCbrmexBdVeBnZX3LH+SnJbsPFJ9sLTuQzGqwx9
uENbw3e1A0ihivBAlmf3VBRjreoG/rgqHl4kzeWC3sIDo5cbBmKoqSyP4OuvzJyO
OYuYwgWExvCTrNK627NNjdj5CGaihQAFR9A2pWbAZMLauQ0uvfIIRd2YH0KKm8TV
RSuKAGu4k+xQ1jeV8M2CjeJ0Ds3EQqFmBR8MrYT4swM107LO2ro7htfIKxc9jdiQ
N3/43wHnG+LXhRdjczfFggBg9r3YtgpSuPi7jmcvnZdajuN3HC3RGzYWDTzvzqpt
hF0K8BM2EqyWlQRXc04gJy1tLku4HZnxKB/t6wMzhUn/iX0O/NN0y07kIR/MwytE
YuLcRD5eOLYWMKO4l1mps4xY/3ezhqNcHMOqcBiK00wc5q1gBWpYqkdcxp3EH61j
8vdNVDiCgD03Xs5h6Ns17UB0RhJz0BY213gfVIz9NRY3YBYAJz4iySw8ThXdJv/Z
VNR+e9qS/ijMzMH+vu3GHY1iddUzGF5ncxJHZ74G3DmlkOhEikyXBsKPctLK1o6U
FA+21nl750WQqJA+spyyf7nwNMxhqvVSY8rGC0ML57wdaAUZPl6eyNf8GtY5ukmg
AakNr8IzPDJfzFoJzGiOqncW54zaEFRE2qWWxrovFFkuLIkoqXEmNR+E39eO5Ojh
mO9DS164nAhWPERs1RCJLqRRov107LgcI25UD3Am9SViPrCTrWwVz+L82CXj7tgb
49idB8T4brT2umLRBsdyvfjnksy+AhakOI8AAmuw7GDl3j5f2kl3odleil1W+ayi
zDFn8ByT0koB6Db0fAwnayPy7HUtxVeYW+VRvOuXlCZdWpcxJQmVpzlbLxZ1ac3i
XD2TNsAc6nFoBvmEbDruDMJMcOotyKeNtku2xsklJmr97LrTYAdDGy8yUYUOt/wX
GNL9rkFFAtSXuH4cE4W9ZSN59OuFydF32X87oYNvgfyWdBI2pOce5ql51hBP13uq
+S6LKlii+g88Xk9BOpestX+uJ3VCIJKP26lkJb30Nj5W3bKxKiCF+yWLh9rthfx5
hUHSCiX1Q6VY8WM+Ls03EGtSMUqFuOrBGr+y0daF/hsckilEMv/jYtfeWwU/iJCs
8F/TE/brUVfIlP6l2ZN9S+SXDCk5WjiPInyRa4BLXgyo0PyeLcuXrpqURMYIZO7j
EwAVcq5TZQYpbtEhS9hEZl5gR2E02YBnkC01zZJR3bfNfCOe89Ls0kmTfs29qX2G
y+IjTG9TLaFC+Qg469CbEdWfNvTjr3c1jgZhLbRylolMMFucXHF2+hlb071Kp/cr
qYpEgZZdS/CU4NjFnO/vEGEWYvApOx7gAWuEYsuU2w2hsuSyTxMkPDeHz05tdl5L
2yyaqNzN3p3lXxnCnCUy0glEMjjL7mA7JdlZIdPF1NFERjweGX/nhHlmCYw1ddGZ
fopmtc3jZlf+tqj2WujRc9cxxjCp771V0GVaA94pi20foSoHydHpPqhYaCVhUCpb
bIP/M35vEuw/Wev0EFnjtQL9uZShKBbwYs6wjWjv7LhEm0lypj8Ssp+4YdwaAPyF
cyMb/6D4gi5OZCrUvwTu4TpNs9oELoOaHaxR8iYD/CyfOKAkxyIz7FhDZdKiNXEp
H7SdHkZQgNYDjCr3wKL1oGzKhfO/zSvxT/J15Eb70VIsWcjs8BvOCT6HkeNGouEj
qt2kujnCvGZ3hham6pggmlnfebX0bFmDRnGuKS+wW2/lXFhfHBxNzy/+d5AUxQ0a
o54w8cfez5EbTzbCljHtYWIcy/Ad0k6BkMEzw098bDJtrNypbrAlAD7luY5kJxtc
vqXu0ks8axsyDfm6CP8a9h8kxX+JuPbcv/mMGy4xavxvUL896IfqH2UHV7cPA3bq
vYJwbt4Q79a6VbyXcQundNCQKz/0lMlTczgSfFksTq7P5nCL+eXs1yeQ5zNPHEt2
M+dLGUdU/pn/eea3dPbuaRBqUbgKf0mrye/MtvBk0JKhOO0h393/YObP220Myr13
xPfmL//q+wPScmLgBMe3+LPIoC02QpPxPWNh8omaX+ZgvKYAzjSBqrGHXMvkYNzy
2u0hH7laPc6c2emg6c0Ec9XDPKENuDuwPFF1kY+FgQ2fXUqYmwMd1N8s+LqysjHl
sOr1T0YNCXOqC7TD4f37ElUKPv9JydWfqVxyOruLhZ95n294Esa5zas4cUfSHXbp
fdaPEFJyr0fMUw7D2ZDeI6YapAYimYbr1t0VC2lEGu9g68sU1z/C2rRcLao4hO26
OnZ6GXRhr7H2YkWwuVez005Kl3l4MUEhywX4EnEwje8JDPR3/e4WO+WIlLg/cBAy
A0CAVVXOn29kBHcok2sY+oSNloxIbFkFo1BclRbV7KiEQXko+nSwxIy4mTWBO2Nt
LS/XfuOZzGoPzZteIEwVEliR313WQ7ZxFRSBvTjifEQZ50PdhA77jLq8F91nFBAQ
Cn8vxnb1+ovrAB36zHRNOJYf8C7wGGzVhyFmoorFeU3mqjGA+OqLXGq+bPcQQMol
WJ84NXDjgWh77AVZIUqBeJlQPMDWeEhRHuVYA6h2nfa9eSCqjCVG0ny1WWnEO7ox
dbgiR9GlR827w3c5Z9HeDJ3WiizGHrDRLS8TTyJ8B6r05DfRmaZv5GjHGDYsZ8TA
Y+IxFIpcx5Esr3+gvrMIwixELGe8yLFijD6/E174hxPK+D694uYcnWvJifU0nQF2
kpS5ZHo6YUx4wyn5hTKufy+dKGzAYvYzb0w3bWNH9ldwbiIcLwQkcf4Poa9xdNop
PY5EZGEsdRWIaE25vpPK+XDLZdqw0EielH+bVDAe4TQ5XEvMV2H3NczWPV16TuzT
ilYi1bwTmXf815r8qU9Jq/3BsD6pEpnCkj5TXQqzIbF9xePV4rpxq8/n+/55tbRh
+1eXq+i08+lza/vrl8hgnmlKvsBOu4SUcVrjyK6JEwTJ7C7RrQhxt47AJSIoHygs
k5SlFHM6vIwiJcJ+ww7aw0aczXvoDDs3yrgiyhOkSpvp1itpLOTOJUCVOlntXKf4
hb+Kyav+gXctmKd1nAPSbYKRCRZUAhHkIpfkJEBytCTpc1p2lSvqgezOGySE8/Vq
aQ7jZ8vvSQ+xusZh/mA9x0E5GirXZb+qJUwqJ+CW+WoLNkZCKKYbjdLxDZ1B4l/x
DtgTyLufrFIL4zxhcZrvdP7MbJw2jnVAcmGciz1E0Zx4X7THc2TYdvpRXLXcdqhO
ubK60jZZFujtNhIzlYxohlmxBLTRmygTnYqdXhXdcOCnVM8FDCmofBH0v1sLKo1U
rlWnYrlHObtvAYYNHb9lImKgEtyUQZceeTN5/1lGrbT29j8TroIUtIdV6nMDrakb
BOs2Tcy2fVwvofJYafLQg/Pdz2EbYzEOn1zINfn9zQbE0Y3qJo6Z90GLnuNHNNTm
coOBb7V/zCU6ilStRGGwOCxYuV+Uare+PSARXW5IeKUQzPD+Q2nvK46GDwsWHsLg
UTaQUUW88ezrcI4WQpS6ncCeo1YVG8Kejh1+WbcWCQDsH2gWgx6VXw9LOjRIl7rj
Rjz1hBdvghpzCrdDyDgIKWij6UNkEA6bMoWwd3GijQZ1EgtnGk3rnqf6u74ZBYTN
x9vdVXzgkQbbxM/macYy7H02OnaYosVqKZ/aIrunCB3Sk7IWT2NLuavsGzDm7XZE
FLRL7tYnrp8FWfFg+n0hflLfNREewGrlwqt5KJBg+1Hvu80CKSiYS7O+LY3juZPG
VVnnXRxMAnriYLsYJMaCgIMKpiWO7KBzUCpO4rVhAPw7byt5VgdztgIdUlkhkMnP
UY4eBSiJ2LaBMaQBhKqaw3mjakmdrUhCTLVYt4BROMvGnP4rIu/rkNGTb8HxKpwx
SuThphDHJ0J4mHyGe9Yvp5lyvoUn6MK06+1rYhkAjQ9SiAHq8O5fn/F3QkYSb0pk
wtUmNxdiZ2b8XGABL3G/Ezol+h7Ess//11rPzMXrglhidV/eqQqMoOEIypT/YUpa
baURjqIrnnGpupjD/tZSMwO2aEM0gu+fe0jvX2eLazN/GwIWXrOrPoghFvFwfwH2
uiImWG2HO94NA1uRN8os/ZRK6ZsKp6VzugQvx6rBlxrD1OZAuzoH2g7wxvoMLQdn
tthUJ6x3t7iGhsIZB04aNCxhq+shRVi8FLlEcKZ1dGKyiwYNwxnPCcPUyJdSEb5C
JgsAarz63Qgn1r78CRo9N/VOoTzz8c8KERs3si4qsXeqFv6RCjc+QGwOkU/+yIIh
TUCxTkEBazSXysz27YA3jD0pnQtK7xvhChpFSv+k3DYbHqrm15xxJOqP00s4lDft
2eh2tq5zshToJ5Yn4pKBV4rzTUFu+TOabii7387IAzcuDeW9kXkblOck7S37G9gx
GtXwEPPN21DXUIBlnHgLIZs8cSab65NVHacH0MZgcRaSsTAtlW45CO99wS8ix5MJ
zD5w58ooj+0H1VtXQpzrtQOx9jjAvq9XQr2P94HFUzaBIelz9OPGlNZgUH8dIrK5
kv1tGqItD6z4EvG2GSlwyREUkkoduFr76i0ylDI+JJNQha6twZcfMBlogrCZQfz5
YDeKYY5y6CfyV6dQAVgONZkHMrcNFYT0tmjPKGX1psvmjVkjCsMg33YM/7JqcfFR
JFZ3TTX4h2Lnhupi3NHIORSNcEeveysHk0mYTcJlg3ofdufrpw3QhPygaWzoUFHv
byAWokIy3PFRCzudzBLQzgHuVC+oWl532v2JX9bthscJEj3iafrXz6Y/JSuhqgRw
Ifx05csMLz2dY4yocYj9sy7T6i28vDDPVPX4xkfYUeeJnDpxTBZn3thkLDbbV4/O
cnpZb4ALK5JSxFcCnwZR3hhmqexND2DB8BH/IQkdpCOgLoHS8yluDzABNg71bJf6
c+va+PhPzxBHmqv5fL5aGcSKpjBLFwF7J4Q6jMHFw91nfRStRYXedZkryT6wFNpL
PNP+HKxSK8PJs8i1U49jQwPyqcKg5FIP1KOl1LA7RT3+kbjMc31td6mNjOBaWMhj
0vnyiNRhffejgsLkeV25Gwrj78pkmZRPpYst9mTEPwRTtAmcLsTSg/+Aw9a6osS/
QY2vprsu7aEzW8BjrT3lOKwFrAVWMygxsHmUpIncexRJYcfA0Uz3iC+mIyrNIrH4
vA1E6EgtzHym1SNsyzsSpieK/PpsaBmztr7jO7hZp2r04t0tfhb+KkAHX/0J2cMB
kWwHKJrHm94BSPY2/wPNVWWVv/yBI60Cs2OM9rSEKB3tgrUoHhqDbZFNPxKRQEpW
QmtDonRqUBGaH2bnnrW/UtCFGEpv0qFb2Nx6nn2qeFRqIyAkOtoGAB5d8sly1cG6
p/zM56bLyMgTt+XKceymuV3krDdDG7c4ELwXg28TB8KWQcIRDSvOLtfbqfHtosKl
450Z4van7OyQ8D39J+AG+LF2Xw8mSFt3q7PbSV9q9fZK3b8Cnr2oCKfpmcdsZ3kz
SohXp9TeEzdLQvaMJtU/HBbNRFrRut/PMmYpz67lBV6WnuGRepdKhXYWzIk1UT2e
l5Zp70xRnnRENKYEB6L1rATmJ07lEauuoH9gL6Ll6cBkj7BiweIsaCUGJaUtjtSn
I3C/Cd4G5vHMTuQ8pXZh3xeN6JKIOs3R+fJv2QC1li0U02Mt94KdY1OBajn/m09l
DSLUnQlB2kGy0/okJeDhPL9lmdxztG2bxb5vw/GP7k7uNo7GItdmrNH3hd8dVkPm
wvEhAfdPImcVLii+0t9kYKXvbLUH4uSZcsHOWt9l6iYwAEHYI5EpNt5ha90NXNdK
fyDRwN6627ZW3wFE58HqfSSssM2MAfcQoziwMBjbo+YaK8i0br+kV2/c+uebMD+g
BGdHhEs5H4woMGknsadUH9WX0asAjeVMU7TyyBLyexaf/pGJPYC+CFAVlOvCpPmE
o9IAfmkarqwAzm/266jivU26Y2orvrhOG/t5y84pi68+mmy2cQGRsLMj0XhBsORF
FRYoAPAopTFTDwrQXD3tYIJ6OlUG2bUeF0zhqfKdrbE4GNSjb1bXxx/uV0hmrnHs
3UY8KHv4Gat1RIA2ZhadI9pY8RFSE7JAB+yWxttlWXuD18fRdpmQtjN1UpGMXQtE
Jpq4R7SeR7RO88n3+8lOnlL9eftbrnjfSjmxc8Zx8/SMMufI0Ornb2zgBaXc4jwx
7gm2oGFEaSxWoWjyiEnjCtifT079Shl0XJtkAPEcF6EFvaav5FYN6haK79ZncVFv
Jpk4ZaLw/hy/JRTqTCIzALet4qpg49KoG2qQ2udEg9kK9GZgXecEYFADLwvXCfcC
dF72NHhcX+L2EyoDHouEX6rapnFeY2RlBl+XkpS5s0xmGXKfVyre6tNNIqiY4bpn
MugJIVZHyNhb7gOZlLXH2DdjTBgP4dmrJxCfAKZsyhEdmPXaeh/wPEVlGSgi+co7
o2VYy3q/+HOav6RnWGDuzlaI+uQ6Cz0b4ig/T6/sZbXpYIJrxFYviWQ6QrVlLSw9
58SlXBkf66csGJDA5MojBea+q6Z5WR1bXMZSAIDRSz2NAsOF7IMiCYbOhGXw9ejt
YDamh2nCkUQckYqNemLHtq6gSB60yX4hJ0Pis5elcML5S7D0QrziH36RLPt187+J
6tPZs9xti8DaTXonL2TBbW0KCt9+E7tZDLMQUjFqYEtqecyg1plTGvfndneL+XeJ
oImYIKdHTSqGROX3H11JZXgaSIhTSm3FeXlVimKNmBSRfR6sxRdYyRTRGwly7R0M
v8cqH3BxQS5AB6IzEoEn9r0AkhrN+Eq8t+X4AIhi5/Gf7NRNN0Qv4Kb9LdehyX1R
R4MJH+VBGPOfI7lqFjcIgA1NDZJF3/o9KzVpu5XwVx5zrze/YWGjlqCNbAM37kni
NhHK93Oo5aEbv1ZJeXYqK5vk93gXu/oWmI+LNT7fxF/PJ7YN/ZbmO7xcllZtge1n
o3H0/Bqu78cCrpefaZj6tVaaiwlHVUFOCwOXgiL4ovfc53WyZxeVFMBR6h3ST4hl
cKCOW4HtOK6L/zxtJ1J2q5hE4IL5EjKfTI+tKbLqFdjoh0pqa7ZIhWko06vVMoxS
/EFEJ4Fb2IOBPt6U3Kg8+lvHOEpGkr/ZrfoP9Cz5ZqxONFM0CPPedl0fU5BArXWh
uM/o+M2FKtwJz3sJmzso4ZMapOF3aql4lIK+rcMiVHDjN8t+IdjPfmuBVRbpDtwH
PYiPEglIyCxlixC5VwS932uUpT2cPnJeZUK6KEK53fLZFdkg6KT7BYLm/EBX5LD3
6QbwDKk09K7EyT5owy8/il6p6flm0K6rgOSzz2oeAmhaRz2KQlbXAu5W2XggU1M6
f0ltGyBP15puhQqwf7DP4gtpSz4wA+RV32tjTBiNdct6vwKHfhybfHTP2vIw7eCN
vFu/1azhStDXMVkSqnuAONmjkDcQek2UD/1Zei0t9ZGcaXy2Mw99wdAhpv1AUk+N
S/D8X8u4T5LSLY5SYx+atzA/2/J/JtyQWaILUC8hRbsg1Hx6bJmJOu4zhNqbasi6
znRmq+nFoHZ0DI1QXRYrg9Z7R4i/lFFIHsCE7vfnHcQYKR1ZdZUGVcBuOefGpV3V
NwPAJ6L+zHF2fuqBQMUHZh6SzWoFqhQW6QFOSjkl3DKpzZ/kgnA+UKaY/qTXnyMK
kiqd2vYSWB5+rNMzaYi7KqxDxJ1PtGqBmmLn1GC+WKXAR+Jkpdpp6CQ9pkgPgz22
4eidMV2j75+V6A14i8Z73gGhV8Uc/d7MyZCQ5/KSKaYa4+1GyCJYpgVtshFLPz03
u5UP4hE7kt/K2iLvRFy1VXWcM5m7zBcbqpARWhOFcsedLxB2GWrdpv3hkAFr9IQX
I9moHBJrDPnZnS7e5KUeilCxMXCNMe68KNlkmOIMsjlWTyFSNl1j7MwRrZaforZE
8E575wENL1SXhqv+Blsf2PBJ3VOqArGp1LPCxTZ7bXtSie1jY9oe0diWPwAhGech
yAwZ8B/Cte0/YEXB5AWqz4rqh/MraJmXi/OKyT/eV2fr1BgqOec2VDUBNF35sv/Y
J3x/Ia9Nx95uXw/NgVsjJohl/CpFqt9Xc95Gb0YhnXmWoH8l9+fOPGwsy3WI1+BD
HNEeXPyaKabP7/Fma3fJXNKDsgX+uls5c/Mvo4ZiGDcIvLrimVh9McaNfgvcZdpl
zvW27GUnQF6ahzngrHUAbP8F+3e0dok1CLo6QA6BsXC2+x/tSo3Gbx1vHYOLZH1l
W1kC/wLl/I5eZEN4sLYOntjcTbjyLL2GgRiHvJ2mcHN/yS5qzEqnLv5ydCOzuCHu
VXoLDE3of/IYPTQ84/pSrjkjA3g/ItZFxx2V62xuFj9ByuYdSQMJcocCjZv8bJw4
ISVT29OuPbkz6dNp86f/J+wZo4wNoSuwE2PnGN+6i9KVMPo8f+y3nZSmgl1b+cdb
M9IwMuN49Yb40iql4m7+Ic2t5vOn8odLFxaNkyXohLLxnf/IjyP9ObSBUDQKUnpc
Q2KUdr6u/nsZW7F46TMZmYovwwXVwvswiAo9e+lG1bfulbmVCorwxeB93U3oza7z
47Ys+DTIcliT3yPUITQm6b6us6RhMQoWJLeI7ghYq0u4de4WVcGmcT0Bj4CJc+uZ
UfPIexOXP3ZFZjQoHEanxcIMJNn6noLo1nLiy4Kaq35UpGr+7Bd4uyKYl/pvaWSB
Mh9mr5oK3bM6/YvYTE1Irtvi3hNnQttTrQ3kg1q4VFW0KTmb+opeexCbFY2RSusU
elAry07peSCRLxoKIghgup3MaNV4FEbj/wQDDuEZmj5anYT58CC1oHXNPwn4GcgH
AVnqiS0g/26CWwitcb2LOODv/iQ6PKvA7+Ihib9yKViFITgegj9E2hj+wlkr10At
HSaQHQazajJhRKl1hNtIm9+EBSrwLZsPBu+3e5BVPk3bRaOWNNLxQ0itIhIZ+k+L
/pa3V7c+G+wxemxWuqbFCs+1fDimXRo/x65PN1ePSijbjMK4IaQjd9s+Qc4r6eJ/
sZzFc+zcbdf7sZcjvSbBMWJymt976RdefIDMlSvej5Knfhq32Bfq5OByJaE0jGXK
UhWLRJr0yDh5SKYuKXqvmlSa29jxbW9H6bFfWkiB/mKGY6TfhHZfQ7w4CR1nNfXY
qOEkGMdz55Qz0mH2KU1Wqb+ZCIPXhswX87zCtKKYTLttjuDP/cgBNBdqs7p3QU+8
jOFUsHPxatxAC3wT7cPN0kWCCwojhmYhJGeEFGt3fdd+Pc2/hZfsyQkjjwd4YB/n
RwuxJJ0i+2Ir9rtb2+n2gDR1aVWBeavZRJnOmF3TCRv3TFgD1qOr+rPx6+/MKG1K
bknDbKQo/m0CfWSX7uF1mwJx2Ae3PurZqw+A1gKqOqo57uPG6F/2B0dWBNerPht6
FONvdb/4ElzbKFh7ZwwLHgkiT1E5+GVLPHxeNfmOktoRwXcofPQkJtEZ5RJY0yGg
nKrlpbdi4FtjnVShJt0OOBR+T5LTJ6XK1KN5zvGIFxD99ZpESWT+xqmSXSagT6vq
HWSlAPZvhqaOht0utkw5t7C5dQiR18SNLCqjvlR5HDFoSTe/m6iyqK4Nv6N2f8/x
XUwvKb3ChorbY3i1lSZLuYSoiMybHx3UZngFq2klltz6wIwUp1f1dknOWnA3yXXb
2CAkykPZGyp7LPQpRH+MzyN6M0JmPTslLoToeYzfLh0VRshU2ey5CZUUdXpDf4a1
1VAfGhEedxR5/hZscNX+bxHcqkIbITEkAbhv/pZPrb0FLu6ld4BWt5WUX8xqZlYd
Q1/hjvlPMVdiKfCATCCmEpKDrBE5lysSfOVEawpjRxyIiGNibB1sPxAsH9wbb4fk
XC8f50WprELdXMwiFFbrRrhWchx5+Dx2qreDDeZn3Lib+NtQBkCM2LXaPWDJZaT1
45AxqSJhXIxFNQk/Vj7KAuDKOOH1e27c1MoaL9Lu5WlRIqCPRFoOnwZlKp603dB7
N+DqQ8U9lIXjYEOnguGiEONlIE2+SZ4cPQnXyadvg5ITYCYuIZRAJy86dBNYF6HZ
0zXvpKJqAlnc71UfaxofY6NDg+AQEdI3XdCzthEzktF0gE6vSoAUIn4pXIenp9E8
iIq+MScaJxfMcymdMyxnU/BxXdcBiIawLal4wvb+3ykpsKdwKsOhNDQyNEr8fog7
aWkNrH/inbkdmnmqz49sGY5xPzF4O80avWM2IHh+aHig+jbeRWstW1Y/wJMfB4GF
Tv1uN/HIzOORaHPzVy55s0CnUnu9V6xO9VcyyyKg2hLgbcB900D9dekKWc/P1jQQ
og4jAmGZdhXyK6RG7GpUV6MPzuH61bkRzY3nbSyK4tMSJBMtrRJByaRniPr7Wko4
aCehSJgAoBAFEbJ2IWXVLBHB3wAUwYmYkYKIEqnD6rvI+XTvaP0obCdczw8C1iYS
puhswZyjOYJCqCKO0/4VvU/vU2wqfd7Xx0cj9jBC6Y7khSkNo7pGGAL3MHp+KqJZ
9OsrH4UrQB+ru/T5zO70J8hZq1dP4jeqsxfFvLyr8uJnIA8Cv6sj9Hr7dq2C2BsH
QHqWgmUPwTaX4+R7MjOIVmnEF1vi7o1taIZuPHmVoyRP7aJ5rK1Y+Tta1HN03uxN
Dy5J85IZaS8hnX2a5lGUUucyYqq+Jiew+mMQ05sppsRx3mJCFzioKRU06sPW8R1t
Zmiywsr9LOdhZezGoA0APlAWRSyafJvJPUgadJtA0pfRmYVzfZNQ+1mOl/F7AGxa
BH201UWiMP2gZbBLXn8534I7CXHNfZgrs9gwmHfiixjBGpASP3KYFgbWOfYWjjoX
5ZKgOiooyJG6mtqzHWmoFdLrlJL/NdSsJEb83mHyZWPNZtoZKF+datTdhjP3cTiP
G6SiNgU/BsI/EtahXkpc9n4FTjbrJKNsICIyLtV3YhwtomkzY90g9Zb+AgJ1DAhn
Q11cgsCAPTnSFZa/dEBDuCRIOoAAr7JZoDMZCIhb0ZZh9YtiCvLoxd+OpJNj/noK
gdLC97IHDmA3j5A2Q8hX7mBOOz3lR/HO59sA/F9MHJe4kHs8NoN9SvZhKCdY99xu
aBOSA7c7VWqiTESrmD4sLeC3byyPHoMcV6mFmzmvz/ZGKkijBJOAYy/1SWMqPzJP
tIj0e8OF1TgGKi/U4b6pk1tvQUTDy5vc6O7iFCRmko51zWNnsdI+ZY6XbIsEp5hD
pTrCV374kItoZ6Xu4U0CZmNxPBXKKlzghzwcHbKYaUbm9fxhaycwLReFafVl6I3Z
ZuM+Iy5k3TEWPrCtadANsqnA/jM5qgxjV48gsFfwRs0Wb2er6XJnO8JOozJQXR9h
DCGOMyZ1ipYMwnbdvTgpEK+sykjsrvPxYo3IpWM4YPNFXBS5qy0TZRDFKojKIjhg
qUJZ71v4YBh4pei91oAMjTfnIySMG2kL81bzuAAqTdYa74gfm73L4zlpyucmzoQH
/lhz42N9j8BeJbpiippO1HxMCcj9eFof1VdlsMHTa/wfenTvqUyrwP2YrZwfg0li
j8mssZeQYcAecuBhZbnlG6MMkhDtDYin/FFKm1UW6bG/oiFkpUeGckF9XRi9TYok
5AjHfefVO5G8/+8AHT2kWr5kUT0/YKp7OVMjd8ebrZiBwjV7dboLi28691KEoHi7
ScPPlBs3vJWypc5ZHMiPD7bBx3lEcDD1DW+2d+ADp1U0o5VSHsgG1SLV8LhXqVhc
Sm0AeID8pRBrxeg29XEoY0RKYKVyp0S/euhPKGsW5kLLsVpnWaxFhmUQc5k/btoo
87Nz789LDsIA6HSIknif49HG0Mtte8OBFpprFvODz7srH05ih0qIclyvhWllap/3
RGa89DsydXZiaaoxzGOa3lnUBQ+9as/ksP4M9SWMnd4RmpakaoLXDVgDgZoSM2HY
IM9qTsLIfP7cBpdjzwKHlOyVa6ZlRVA4gPwJix4MzKEFoxKkQjtwbR+mr5dOJ+UO
N9whqsHhRGTF1dxnoTCn1xfxMdHM8UoX2w77z/jV1oHMZkCTJYx/KEQ7Fhv5C3lo
9q38znxoRzY0dxUSE7SFFz0reuCKZy3LyfgFgXIN7dnjWrQ9OzTeNYgq/DcGz8R5
WATNhdOVAX6fujxrLncYCd2/+h26ipV5AMTcGkKxK3BWB3k0Vx9rZmVebYt0hVs6
rR7FXMhSFgoVfdr2D4GdKEhdWU51441oMgBkFqt1/JgFzyL5b3gMB8qmkZeTSNwa
ywBsB4q/Bu6Q/4afcZff93EiueQ6bJask6EoTBWrOiQ2gXMQ7fr21yI5HBscmhIL
QRwsr5u08MXKogb4D2jU7+w9NUSBi17bI2e2cIKn36rDak5XsmCKs146FMYfUg25
SEwjJ7Z6EPq0/rv4GLNLBjxiBJocrmFQHqHdzZRpa31CDzy3X0hjGHZZzxQvn0xn
khrISOIFr/t1+3hot5jB0UuEPYvd2tQZWSIxVbeSRRZjpNSynlYB1hD8/1qHI145
2oAC+XfLHTiXjNk9NIOszkSilRzFG5IIh7lvXEMNw7DVFiPYrhD27rC/uLHmRIqC
R+850paVy5gMZ6ixk5CIrWQE6keeyijkkM5+Dbgp8WPCopVxywEm7mqCzOzK6hUx
4wp8teMWV4xTS1dkQNLk1dDcDc/necUSO6Q5HYhH0BjQ5BMwv/IB/9QsKCwI0PnQ
+n+DcFX+IXsEjPYl6Bwa17QMZuaWOzyrIresj+OB5Mw1uh+zu9umDyZxxa6VBYL3
gHpgYHwaKOFhMhqvpe3rcqixv6/YItid8LZIJ5O2C3w88VM2Lgrhp8TM7dTEWzB5
0U36qaeYcFmCDQRFndqvOeH4zt45d1Rx1ACd50nJ6ifckCt2rHSpFRtS0+emqfhp
BwHiEFh7KHOMpso8JIIh4yOzz4/Vee88ppHkiQ2otUjFriMaAXlqw8Mw2u4k1p6r
PQcbIQDqeA6BteKO7pjT6K28vWNlPJOWSBJgxtdPgK1AJFxeZ6j/d7vh/rvtzMBE
jP4S7oCKizb0S/MpSqmNsHq/bw36tODc2ChxdAMXtqEgBIJDHVd1g3N6W3/UnAlv
1vxhYeWDOMmzW3CdD5OhgghCToh46jN5bq3jpXgThzeIfm+XifHsdQf4Z1xU77Cw
bj3E8V1RwzPULq9A2AEYVkKBnbe7FEKYXMPTV9HQPYnm81Hbtzoa0uYRusFXb/O/
aXJ84va5nErIuw1hg06DKJ96sqlqFmJTK64bbc6M2tCQKzpq+iaU23RZcNVqRNs7
jOazqwLGsrjkXTeUssGhezMnb7YmuhA2hMcMtNgwZAWjI0LoE/Z4fOnbxTAGaIUh
MeM2gxO/4lxB710JfygnONBDh8oaa2q347Uvh42i/MvlNuZUd5LDw2TEssBsSwj8
gwq2rK/IuL2tHQwYHVeB3b42QkotuGcOw5nCZGl2pHovVGL7ATTK2dUFKyhZe0oK
gC7VVRCE9tTL9icCioFfEOIOKBhqiyrDME3KvWxznnRsa+KIid6Kfekctmuzh7a0
omezqy5FXsO8nD29AsC9ThV1YAMOYwFf3AIapilgQGDA8dSqmieJgCKY4+j0EmEa
ay9wOfPI1el/OwJtsj4+YfQfUwaFwLiiYmq6EdI8MjD4UEFv2e2D86hCG3jkWpKb
DClr/caDd9WaghL4VvMO5Y/YTsQNCBghthb7VjwgiKeX1J4hGZAQb9zFcbHQCvYB
4bSy3Fa1M1//gOBOMTikZDNXN/pGV/M9LZCtNiRppSn7O3Kelm06EF2hdEeor/KL
oCJMq9667Z2XplAloD8UC5T4tOA5uKt8SOTq3n08wHGTkVtn8gdu/xV7q36mMhFK
UgQdoT8hx4YMmicLLKtfqSmr1bRUEyauE1XVuUsd39xXnV1+5ybPh8fmCxHgJ/8t
JveuP3HU64y4G35nfwJHX4AKn4FPiWwKDsFVy4mHOvVys+il8lmiyEZ2WVVivokN
b/f10oFdiOOa4OpO3mBgwxMampxJF8lQPM+Eebic3bQVx7cuAEip0YOC/xxEsBMx
3agzuAOiZzOs8z+NLwAc+0F2fFWfMIXCuWFFxaMxtqDbycI4H5V0CAN0WXv43qo1
LZRKDxV1LzQSUpVcefhPE4W2b63MSTbQtjzIw3DJ1I7WEd2hblTLbT8XlCWrVpwc
zQyuQcYIKZyu1xpjoV+gESjVlD+wWnrAmrnyUDhu8LgUqfwQwsUWISuY9D3IdpXT
HYDBfwcS1zglrW+FKT25tpBxfmXRW18g4TGmc/WH1OKBcfs1OiCakoMcNBA1HR5F
4AiSlb5mq7IBvT+ztMPJZLhv3wDZGPV2yJWVtqygqU/6jCDIlEanFKXD7oWUd0Nx
nGrvUHRTGlzWdCIXOz/EISGwO0yngBKpESLq/XrkIDp2fEF4YNTGJ46devZjlcgq
E9AG5kbVqZ51HdQQEH9CbZaZa/3Ob02XLf8ECc6sAka5THemVEfAjOqbT7KN9469
BxfpEDGslDcGJjkQac2mBGOfV/37bBdMufutBF5R1a0n9m4cv47bDOr86C0esjjL
BUHI6zN56cCMplxNlzSGZTh1ILE/NTHtpb5wNQ9DcnR4vTdMUl3ybfkT5u8SKJZA
mORl4ng8RF2vMspfE7htvGZGWtO93Kqj+TCp5DkGki5L67/jM6RRqIdhMVwX9EMI
oahvigsBjzYBZgK2tah/b3M+v/h9lg4rO5U1WLOLsn+fz9FE9unJwc3RVdsNsvbS
tQEuRQJkCyF4/hUJVf7KoEBf4TuzFge1gqlYFs8LJlvzSToQ0z1HE5FjA+lqP40e
fsbZjLfrtxAyxWL0D6E3zZ3KQWopQxSjWm2JBSrAQ7uqNL/a4AxV+itl+/hiAald
sAJxUh6cxj/X3GalGQc4yMU5VqL0iVLHhGF9BV5+IoDreZBV6LnGatsapFtA0Ej3
cQ6UolryD7ezU+CKiBZR5rgKnMfZd/LnaVGlZAso25E9Etq6NOkrSUNpjDISuXnU
9aQMhzJAnKgl0+hgO0/nmJYXg37jP/OR9hk24qVciNtZuYVJ84EsPUL40jrUQVSN
pPz9A4fMToR0nyrP4JVOCTqaFhE0esvcdaOpRiqKL2YIAMgw63v3qrAi2KwpJwVf
xMpIN4lX/J/3/fhL73kFDkqMo3631EmpVx3Lc7pfji7onHDEVMKfi8OIYoEPWWNW
BJzu0WL3ywhd8fXhg5HnDo7YPyQjyDBjD+hqmQCQSar+lCRnZBO/UdH36CXSmv3F
/i+38X4BJt46QMdZOx/4ST4TgXEf7gwv1sbZaSkXLV0yA2QONexo8QqynY/QgydZ
i5U09nBpL6ay6aXcOdJnoNksjbjoNt++3VlQJBwxqqFCVaw3DDcxnyM2Yr4j1hXL
eYaxj6MgJ9vpPGvSld2+ToSKT0QQ8kkij24C87S0GNCcot5NFE7keuPT9jOa0cLI
lnOenkeDzkSZ+IzefaD4XmaYlLG4Xd0zAGZ+rih+gfEoWhF4DrItTQ88q1sesEgn
wCrucaaZH7MJk2/XEuwqChjZeBdItD8FFRtSX0haJwfkLByhgKtBH/urP4FMJJLX
Ezk3zRPOD03vDhlY36PIV4GI4PXYEQbt1twIXG0pyAJSsYmERayHNwrF1NJ906yi
XN13ccl5hsMYdRcpC6XXD/doOJHOGqVUgxsS9ZMtJWLhocQQdXP2PscMOKLx2Lyy
QYlK43pJoEY+59WvV+MccbIeWeEMfIyvFqtUwvuGrakD+wkDMzxoK9TCjMuYx00Y
WOlsLkwLQERX2l46bWw2tZRO9QF/8BSPDkDYtfq2uJ1S6+LA5XjrHNsqPWuWVU4a
Ch/DX7CuP69bVil0gxC7rIiE35JQO7LHo52hkA2BHbKrtDYs0UysQW0Wf54TVjs7
u2v4OJYOHY0cVp2mwh53kHcc0d9VqqmFNw6fX7ZbleyamG9/QxuDm8/S6npdbXF2
rwhcdDXFBBSRLLF/mDlz0fur6tvfoB0/OwBf80o2JE5UHcwIwsohQ7FOwwgL5Nua
dcHp2oiPgeQUV6hAJCWaHPYIQDOtM6XqSf18fenKCBRevYWzsK51FHUXTLcaDr1C
CENp/sljw26N6sFtbJuNQ5yeSosDjk4u3N96upFuciAPyelHvQasX0o+eH7L9t5j
Dx9+AvwvMz6cXCqVsyEUXi/fMpCa0izLmg0Mr4yQVpsGgJE3WdYe1GqCAkPKNGZ8
pcSRuV+7B0xAvhUiW6AN3CC/y7njxWnSbG8CMVkPGUOpK5eL4QbeBpqAwvgqAmio
AAebTwDy2AoUFlopf+5M8/ry5xTnpC+NJmCGTXUX0/bsoX3O84hEZv9lVvaQFM8n
7X21qFOIWVJYMM6IpaVkZB2Z7FWyZtbfBwqkYKONvmuOnMUC2FlcstRiMF6N6se9
AQcOIE6jEZ+f/E70t69t8GxVV1vwVn5p6yiKirCO5yjNmp34m7P/FDOq63j7rhjX
O3C5rUNc3/X6UCizH6U7drKSWA+71ztMuHQS/58JOCfMVGupBvCgk1sBR4oe8H+D
Bd0mJpUBGMFpmC1qrw5rF5XAfuSll9gkJUZ43X1zs5yjnzZKzaoGKxhAJPRN8h5X
EhJQW58+xq1anrhJkIyng+ZSe/rfwGzrntDxc24yfxsnU3Rik/7z7K3ZEXsWag5P
BwdayveRtruZrGOC0nsWoGsZqyKelqwBxlmuZi7waAgRZ6v+X9s8kP0looc3Z7a2
GP9ntBzOdIt9k9auN/bppaeAOASRm6J7bP/HgUnaWgTfzqwMBkjQdRAjMWwBzxZp
RZfIZdlWvf+MuMLuBHNl44sBFHiGrvkzdEUaFVfYxZ/YXvrAFPhWShoTtiIEkls6
coVblojQRoti3mjlf/reagQcr3cYIP2xGJxH7UsjHptcEnv1bF9Si+AqBvmaOM3n
Sluv8IO+Ee9a9rvTwrKHSqSNtw+mtePIvsCsbD9P6hGtjcnEBrckf9lwL5C6Z3qx
zY30rZZ0DAmrl6eMLvCnmX5yBujVWXQqKPe4jxAdmGSEoI8bGymgp8zK8WAHlxuj
WL3deP4Y9miYo0hPsv2WHxDs2DcQdy08jC78kzECZthU6TuMsPWlUc5wbI0NOvws
FQQfj+XK210B5+P4Jw0EYMa6claN0aWzOvOIRHwBjHKSFLw3he+nv9baPv9IH8yL
HZ7B1EHBRvje6DqQrNJBBhayEnAKi757tFDBFOCWQCHKMIk6BJKCmllvOir56q+n
K9sVaGPXQxSCN7WC65hLyiiPRreQrEGId13qykAROLze7CxybdLXy2sHjA8QMxPM
dSQBGX71vtliVPLKfkjubxPP81vmkg8SSdrW29tUkkcP+BupH1alhBl8f1lP9e9I
8KPfqbni4IiLopY5OLXX0u5RKO769PALbfkhABOWzSkcSa6XXubb/3CwaniS/7es
uxmvFtjef+PO6tBfIDMUwwMoTiOX+kqVDG4UFiQDUQPEO3YBtfBoA+ega34ZNtiv
tapD5CiGXmdptu6p1CDsX/mkajuffG6FPaIdgdPT8RjZe8MZRiO+d4fPCtqoeRlm
iQI56ohxWtLL0NJzPT+oiiYDTSjydjNx1dSXvOpBhGnPbkFugxXOW5syyfmy6q8a
NWXbYYGVsJWdZtNg4Rugpn0a2wlByjxkWIy5BQksKw7DrZ5/60aDG9XQDASYskI8
m/oWfUXsrd56gQTjKGOQrxF9Pp3iVfYFbfSt60hK/onAu3T3NglgegUy66TwT8SF
D970EhpeKLXnqLBCCWrAspdpvYvtSmeiA0OPnlP9qdL7UE8Avo/en8oJvyifzZ5W
X5YZEY4b/Wm84QSkMhSd5WiqYbs2I2dgE3J+/l1c414Tg+7mqVG5UFif4ljD8nTf
+6aUrPpFE1Sx3S1Ih9QrIIP5w1Nxrd81t5bnGZUF7pKa3UDA0xJWTasgPHWwijMU
pwrjhGonubrgEe9RHDxz2k2AqhHgM3/Ae7nU1Cp9DSg9Y/cOw7qXIS9DjvYNkhw8
jroZTH6LpKVi5OLM0179tF2cVWniBsofcIwY0g46WkuYVTQ/SQVyuET2i68frpJd
6WLsWUPGtXWHNoX9ryzm8gG5mwn5EYHRb+XpP1kyEu6gVGYxwM3BM7sZdYE15bhs
LuUppuwN9wGJFqyOdIzG4KGcer9i+i8fNZA59fQHUyNqM8dIIpz+HyR1cHlJuuei
IlrENSIxTiTn3KfR2QsqM1aJd3H82SpqZ05zQp0N4lafU3NIxhjWz+l/PHaXPkJX
8yAoXGFPLsohNdE0VzQHWwHBrNQcp81pCDJgjGdU3J4nxBxIJzmVUR88vhwRHnU+
zii6/9txYg5LzNKpadG+hyxk1gG6gmqwmheCqNWbSNw8+JO2LA+Cfmx78QE3TJUH
i+F4yj0Cp+EFF0zpTJn87h3rt9xtOkqw1GtYkJiNwQWOMw9OtcOW0p7ecAW5AeT8
7wCD5cZFaODj9tJE1BGpJC9+TqU0sELqhJ0401gydf6YQDFaNZ+swf1s+jcIl1+o
m1b8flDFykBwO/r0/5agCiyUtRx+6Ttzda8l3QCYUM0Rig9xnOS7UoHEQOLF/gZ2
wMuPInpZeyMqEW+nz9yjH5tvVhCEsxPR9SRxQ5/+nRjwvg6mMFiXKOVWWx1QwvQ8
dRWsipDvIN1ewXmLmlGwcSrMvdrMMGZSnnyyz5ye8H43bLPdOakLZUWgP+tXLQ2p
TEEhIxpGzPO0qfenUcWXIc7b5RCF44TOzSy0VeudVwLU100YoYHga8uWSe9yIcCV
IbjDWtM25J8rchuN/Ynje//Ycfzx9NmX5i+8AXWm/tFrX6QDmM80svH0Hv46HOST
1zTLo+SAmcdQm4wTxRb4ru22BSHAlHpq9qoiPrt6rkDrA13Sp3D8KgRocQgnoJAE
JALcrAqCtetn0IyJvCozwi6dackEaSKCuFQIdDZmUh7GWF09BYye9ZD1CIu011NT
x0xAGE7Fd5DqmjR/Hn/KF7WO06E4gNN/pYIHeiDjBEmnohFjWL6ZuLXPinz50AWf
ukX4J5priQD49O80GrkKhoX+qVL9fhtW+RGFr+juBlMwxFYSZajzyNUiM8qxTLrg
l3DcSQgANiPXHJLV3GpF+vXutGUcgjgPZQMGO4WzTozSCTr5OsQAlESofjuSmXPW
yIklN4X2C+I18o+9RQfWfBLJkXQrjI7T8mkS6pL4hCOpmKSrkRFCV56vRNMWqld8
o/lV5rSz/bRL5sl/7zRj4ZcMJEghQTnpEmFR0ifM+gW+4Wc18h+1d3N3EZFI6hei
HQ/E/OtOlTv4yUz3aDMbV9GT3EFWNEVufjFyerI159RKrer0rjxt7SjDVHZS8YOt
QwrU9AUXOFk53iAiWj3E5U4r9OrzBkDlu6n7RagzYcyIgU0vO6Fw7iN7ldKmNFN1
TBHHOrvn6MWcuwKxvEbRedXd5M2PwMVPUlix9jvieusHb1oAVrF9sEnTNo2PblUx
VGzzIY/LGmIVfR15miAWWdn2gvTVDQvgU266OAiLzTvYpbmO3iEg1yKO8+nmo/Sv
XsLIPxz3rQUPFy/bL+Uko5J1jROmocmEf4IAfjt88zKITH9oTeFFj1MDQjIUdk+u
ovyZmHnej6KNfqLzxgJK+oukjiUfSofMzxOMSLrSL68KlWD/0bd31AXqD90yOky7
90nAHrgJ87kizmzPR71bRPZUkLMOnF29EEkhqqebOwkR+tVWimM/V96W0LHcD6kN
+cgKVhWjNviBTVaUTzNZn6sldVp7PEm5B2lmcU6N27PrxvBivuoaFq3qz4So2DVe
8Zt6vI00Uy9x9fvOJhRahM4YARFteIXGePFc5OhNY6HkCOHn7NXJ9OTCDEAS/q+R
Pm41eEMG0XqZ6zsK2JeB6+gp57YEDJtM6KjElQXQmm8JkGGGsmPiWS6BaG1Jgtm8
jbZQCw4pYLKxur2adGLuwhTmdg3QtCU/Tx9uZJaDLnSwy29kkvxqYvcuM3WS2b6Z
Dzq9xUme+RWL9KjDIYp9Sn2D9ydvCo0quwMV8VwaOLmhEiTyHbRXPTlxXUunAy8c
439uBy2Ge80KmLQNJXE0FCIYSihArJjVujt8EQkpp1ZzOjCUelVBaJY58agO2yf0
JdXuBMrZYaYxisRfuAvNrCp06LFiyfKDl3ulq3mFId3ipaCLR8sKboA2r/ZK6Ol5
WTsfGj98C745R5ssBpzmf9IFSy7HbeGPcnJUPTituWIHs0YTtFN1s20H5pddX9ut
qgsmAw5DXcajtBJGNmmLkzd2MiBF39CHVLMwWkwQvo+vbZnwiGNyX9RRnNwtAG9q
hN6kzTjPcmN7Wfm1yTEDMTdkGM2Oas/vgC4DrJQU/xFNldiPlThcFiyY55eQzTYV
aVQL2yrLa1OUaZg0P/cwPXqgw+pn0de1bTSeN6ciSxT/X32/VzaN9PYxaLKAyYlR
Vbfv7Yzng3PTa+1EZeI95dTWlyy7w0jR+eS/+sl5pQX8ntzB0iq95ZR2xScJcSCd
R9xHaUoLoVhnkhJJC7b4qioifrEKLiELpWpUIfD38OSf0wjQG98i87gvI9LvyUDl
AsmwklY9WIM0r9m0B6eCwLxwIWQb1LpMN9fAJ7UQDHVwjJ8k4vP1Bg0o4U9Qaa2x
oziAR+Yy2ZF5yRXi4/NBAPsjeBGBs2n2jES3+ym4bZ/8hPHyY1HffML8pkEsQ26P
xOeg/a+ZuzcpQcm3ulytqDk3WqNoTCB/9qCC4EjWyWnUygBjv/P0zW8YShSRtZd7
ayS5QMEB3/QLvHhd/cs8SY2GNMH7j8FX7OV+GOT7d4JCfS4XzLj3IVFaso7YmZLD
4HWu7P3pMPwUripsE4Nk0DdFt40xUXmPG5HIaHpBBVBeYGLebfueAptf42vzpd84
jaJFKeyBHGbE7TT5FREvR8OOjGYR11TSfZatjAGZyd7sgzO8vsWDmspmKdF8cK0R
HbZ4vSbv5/GZg/veuGY4ezuIm+OD1VYVc4wMz3TWQrwYInChOL3i0AvR1qR+9vwR
sC4miBZ/qSznyi7EgN/IIVuet+4Y/7VXasS66pIgB78/NjHYk/k7EcO0WjHCW3KI
NUh5BzKi80/jlKVynPvE5q93T3+ou3eL+YovXqo7RG9TlH5ikeGQuyw4d8weuW94
jhs7PE60zwdQznFEe2jVHOkcGHi94P2kjhP3j3ku7sRuyvUJTEdZRzC9zzf2vMAJ
ggUb6U6H0JSXvjTj5BI0f+i+6q0ighH2f4d6fCAIoKNuI7aoGzzbkAkxvFHBK/5i
wldP64RpTKrdbjaj6m5T9lpuJVF8z/DCow3+4Vczi3iSm+SMGcowTbK5nHc0FyuO
n+QuDE6D1B2CMlcWh3ExLHNUfZv3fdUKVat1cMYDWNTi6jPu8PkQU+SndHrq72Ri
cU3IHj4TjPwkYI+uoJ48tARIl97pjfSeqFzH16nCFtOXIST0vd9cznmPvLJjhlF5
JWo0NxUDARruxK85hQsrrIm5nyxMitg0OqqKgM/gXAMNMqFgAviJVDzcU3S63Qc6
JQ0LtUzNMJPAeDw4xKQXM/4GpvgVBNlOIcTBEK0oxuZNUee2FvnkfCHHq+m1MMIb
RBk/DSGTYffasG5ozNpNu6bmujS3l2mG0Z3fkME16zhZcxxFsD8WxQKpkBqa/Lxf
w6Z3ch61jwUF4MZTzS5P/3CiwRl09dfd1W5QNjQ6vMRz9zZL24RPjOVXicX0fDZO
pOIxjEo58DlYVdBZOyb5+qLz2ntZcE7nx0E/gSwnHzFIXcbVo8Wf1kmB96RwFayV
QcbK81Wx4AmS7rnqEr0GL9+9REVRPdwCpRxkd9cZ96Buo3Zu0cbgmnWIv7CBJewV
DIR/HkVkl5ww2XQLwBHrWdg4WaYZ8vzcCMW/DVzfakXrW5GENcNn+YY9vF51ZD6d
W/NsdHdEtakmztrCv72pZGknkxERB5HhtTElL3nO24i9FmLUyPIqug/CAaGzc6sO
kouEbqALhOFMy7WysXeccQmfLWSx/PmA+Hse7LqcOWwPgu/E1eS/+EuH3SK8APsU
S9F3fT8NlW2cpSEey7FpYNnhsREd073Q6lOT8Dyx9F60zZWaZi4o5uwcZgGlioPj
gu5WHipk2hktM1Tcexcws8not7ET4I5PAnXfWnC6T9srebwsHjpp3zYeb18SOSqO
puec08rcckhazx8Td1wvY1rPIUy83xWYoGsH+/N4BN1ngutWYhxJVoKGQIctG1PW
0bOqS0+lEv+a0vFzvVtQbDtU1sUrsu4Mv+QjlKcBmT9bJU3woheF3BsqOLLVe/IW
iI7hzSQW/xMFq2d0DRkKlKNeVAYHVoDp7PmHnb1vNFuwDiofsecWXkHSa4/etTlg
oaKfgUUPfI+YNrYuMGDvhS94GBJmgn57T0VHR1BSDaBetRYSiTPBYA+idt88G103
NmbcmwR0YvjDCZpmjzq7+EVo/8BlnuiCiwwm5rrpZAbAd1QcVNywuaPSUMjsFnFd
KhyEfizccsTRwE8d7W0tzj0+a32LJsQE01YTrttQ7n17mgQqQrnp2HPJJ7q8R4ji
hPDiBso0W76mkrDAJ1q7RDLPTJmhSRvWOew136D/baSmmR23WvXOEpm6dYrBkEUX
2c9F6xQi0xfC/PdYq1nZ/mF9GPjmyOwbbqwHw+wUVKSH1JCfkLY9+CnhQU6EU4dW
JnaBcNP0zhWCR4D/CMRKZAxQV85loGX0uA4gIUn1H0UJDaLs+BP7HgNe+hJhiTkQ
WXnAl0zx9QcUKyJq7bkEgtJcP8gU8hCmD0MU0v6BwcvV2ooa2AlKpUpqo+XVLFN3
KUvvzMWYjhY+lNbD5M9+BMmjZyaG0J8hrOSE72qVPtNf6lIBdVY2csiQ5eF22GlU
E9dxMSO4bBhNoQeoVOnvGAMpA/haWKvmotplsvOWoDDZ0ZlSN67/c6+bnw9/EuGP
TFc2BMtq8DUiCSrAfdpuOW6KI/6Zf6zdmkMun2dHP5QHN9qQYn+o1UoLxkD8GAZM
gYUtljHOSvk9//HZFwEIljdt7VmQis2f+9Gx6meiKdjB510xbhGiMMXlrpliULxL
Lag2ZRSW+6oecBQw42ig1zUZa+r0v1ZNN/JccRKj141HIeiacgMs15cv+6WMVYbP
xN91VnDcsNVl8oc3XFNT2d4pxObybXWNkLWIqq2OoQ3OYztqDUeGo0TQqlrFSqzd
9nosuMPb721pb23Wz+P+3D1QZNC3QyrfoYvS4Jiq6mZ6NRJnaTuk55WgTbtmYDnl
KJq3QUrhwkst2HcChiOMvHnlSOKJey0H+44oCEhjYx+g+I2QVMKLYwDaXvcAQTuu
pECUokUB9gzau3eof7b+N5xA9bD2JKtCOdpLwZ4c8LXY9JcrOcIOZlSxXyuQ/yz3
f9vxAWoXA1kg0xwPvUKL8U4zG1XNAyAt+SEMX/IKQXGcR3xDa0XW5HRJilozTfct
/JNP6vjOtTwgr01kLZvCpcNKfOuer/aI6HC13fNMlFSRkO3fe7W4jUzoTtDDzIzF
NiHthIaDel4P/zE20/sVHNIwxorIwUuFpcaMcx24EZFxlxY0ZdkiK3fHmGotTzDD
DOQ9dt0eQj1Rrj682DXA2JLbGdzAOGSwvl4AwvOpWg7R7vOjVL+Vz+UIbaXxoLlb
AWzPkdOq5uninCICMnf4iQKl1WiJowsHJYY2qRm5uBQSYudj3xcOvSunKf75jiy1
nIxTe4RHPMUxht/dmM07C0oKL5AI8J6nyfuqyRMhIdtzyD19+79baHK3aNw0B+VM
GTrbTV/7LSwiBaGQM259udex3SIs+JeeDW9Lu5ut4rV8O/eTr2/roD0OldNUKEmu
OIS8OXNHIMhJ08gjBhyZGadfc8j40qJxEHNDRrnRXfREBsRnEBUjWcR2bGV7rfTJ
dgPGaMX4BjNIGw778E8wonr3lA8u4jIdYbCeqeksSO63oDSou5zYayorgbA6gr9M
6/TcPtjShYzDuE7l2b/a25A/Sk6wl5FGE6li5ewQq35DeNWaEi3d4KMsUz9dHc64
K8OmtzVXpNbq2VkRtqWpPc8a3EFFX+2FUbkTTOmMDW36w0B0tVLGK9wl8w8cGYxI
XgoFIVwu6zvTY8rcFWFQuLSV5BYAoyizQ0mncgdCi/A/Pt4ExrSUTpf7SwCiLaxb
bq48LCPE/oYaUmdC+CETMRb+hQoyAVDHpu/KLRQJqUxUYEIW9TupC+FGrVJ77fOi
ZOjp+DW0H4hEQfQrcz5o7/W2fB3bgj7Mox+ZBzLIIdRYgOe7suvPSdtVEQnGtRXT
oYSAjpAS+Fa6QiTs9q/ZAqFia2f4YRmzHvCs43DrfBBwqPnalJxh0IlMOmRTAQ7w
KKJDhMJVCh7I09lq1BsRtVK9K26E4VtSgbODM24nrXdFEl9yDzmfoq827QVD6Wwl
qXyXurXS1osgy5jIjtyKp/cJrS76ib8ZDx8FvPTLnmtFzG2WuYo07saj0PE3uLPW
AZCgvuR9jzbWGU4bxZTteGGMxuVr69y0IOMD8cgHxDzogyGFOGBcJhQgL5/nTe0w
t1lkKxl9trDnfFGN8FHHP35MJkzyYpYkDbTJQHtua5DTMMB9bcyeMl5vIdte3uH2
0WvfE/bAwoQLpp8W8oi05CdLhSmBDQRwW0PMdQQc6aR7uTqWhJHyKQ9GuLJKaCVc
`pragma protect end_protected
