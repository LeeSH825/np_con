-- slave_template.vhd

-- Generated using ACDS version 21.1 842

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity slave_template is
	port (
		clk              : in  std_logic                     := '0';             --       clock_reset.clk
		reset            : in  std_logic                     := '0';             -- clock_reset_reset.reset
		slave_address    : in  std_logic_vector(8 downto 0)  := (others => '0'); --                s0.address
		slave_read       : in  std_logic                     := '0';             --                  .read
		slave_write      : in  std_logic                     := '0';             --                  .write
		slave_readdata   : out std_logic_vector(31 downto 0);                    --                  .readdata
		slave_writedata  : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .writedata
		slave_byteenable : in  std_logic_vector(3 downto 0)  := (others => '0'); --                  .byteenable
		user_dataout_0   : out std_logic_vector(31 downto 0);                    --    user_interface.dataout_0
		user_dataout_1   : out std_logic_vector(31 downto 0);                    --                  .dataout_1
		user_dataout_2   : out std_logic_vector(31 downto 0);                    --                  .dataout_2
		user_dataout_3   : out std_logic_vector(31 downto 0);                    --                  .dataout_3
		user_dataout_4   : out std_logic_vector(31 downto 0);                    --                  .dataout_4
		user_dataout_5   : out std_logic_vector(31 downto 0);                    --                  .dataout_5
		user_dataout_6   : out std_logic_vector(31 downto 0);                    --                  .dataout_6
		user_dataout_7   : out std_logic_vector(31 downto 0);                    --                  .dataout_7
		user_dataout_8   : out std_logic_vector(31 downto 0);                    --                  .dataout_8
		user_dataout_9   : out std_logic_vector(31 downto 0);                    --                  .dataout_9
		user_dataout_10  : out std_logic_vector(31 downto 0);                    --                  .dataout_10
		user_dataout_11  : out std_logic_vector(31 downto 0);                    --                  .dataout_11
		user_dataout_12  : out std_logic_vector(31 downto 0);                    --                  .dataout_12
		user_dataout_13  : out std_logic_vector(31 downto 0);                    --                  .dataout_13
		user_dataout_14  : out std_logic_vector(31 downto 0);                    --                  .dataout_14
		user_dataout_15  : out std_logic_vector(31 downto 0);                    --                  .dataout_15
		user_datain_0    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_0
		user_datain_1    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_1
		user_datain_2    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_2
		user_datain_3    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_3
		user_datain_4    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_4
		user_datain_5    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_5
		user_datain_6    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_6
		user_datain_7    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_7
		user_datain_8    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_8
		user_datain_9    : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_9
		user_datain_10   : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_10
		user_datain_11   : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_11
		user_datain_12   : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_12
		user_datain_13   : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_13
		user_datain_14   : in  std_logic_vector(31 downto 0) := (others => '0'); --                  .datain_14
		user_datain_15   : in  std_logic_vector(31 downto 0) := (others => '0')  --                  .datain_15
	);
end entity slave_template;

architecture rtl of slave_template is
	component slave_template is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			slave_address    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			slave_read       : in  std_logic                     := 'X';             -- read
			slave_write      : in  std_logic                     := 'X';             -- write
			slave_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			slave_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			user_dataout_0   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_1   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_2   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_3   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_4   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_5   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_6   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_7   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_8   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_9   : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_10  : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_11  : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_12  : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_13  : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_14  : out std_logic_vector(31 downto 0);                    -- export
			user_dataout_15  : out std_logic_vector(31 downto 0);                    -- export
			user_datain_0    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_1    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_2    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_3    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_4    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_5    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_6    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_7    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_8    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_9    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_10   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_11   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_12   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_13   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_14   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			user_datain_15   : in  std_logic_vector(31 downto 0) := (others => 'X')  -- export
		);
	end component slave_template;

begin

	slave_template_0 : component slave_template
		port map (
			clk              => clk,              --       clock_reset.clk
			reset            => reset,            -- clock_reset_reset.reset
			slave_address    => slave_address,    --                s0.address
			slave_read       => slave_read,       --                  .read
			slave_write      => slave_write,      --                  .write
			slave_readdata   => slave_readdata,   --                  .readdata
			slave_writedata  => slave_writedata,  --                  .writedata
			slave_byteenable => slave_byteenable, --                  .byteenable
			user_dataout_0   => user_dataout_0,   --    user_interface.export
			user_dataout_1   => user_dataout_1,   --                  .export
			user_dataout_2   => user_dataout_2,   --                  .export
			user_dataout_3   => user_dataout_3,   --                  .export
			user_dataout_4   => user_dataout_4,   --                  .export
			user_dataout_5   => user_dataout_5,   --                  .export
			user_dataout_6   => user_dataout_6,   --                  .export
			user_dataout_7   => user_dataout_7,   --                  .export
			user_dataout_8   => user_dataout_8,   --                  .export
			user_dataout_9   => user_dataout_9,   --                  .export
			user_dataout_10  => user_dataout_10,  --                  .export
			user_dataout_11  => user_dataout_11,  --                  .export
			user_dataout_12  => user_dataout_12,  --                  .export
			user_dataout_13  => user_dataout_13,  --                  .export
			user_dataout_14  => user_dataout_14,  --                  .export
			user_dataout_15  => user_dataout_15,  --                  .export
			user_datain_0    => user_datain_0,    --                  .export
			user_datain_1    => user_datain_1,    --                  .export
			user_datain_2    => user_datain_2,    --                  .export
			user_datain_3    => user_datain_3,    --                  .export
			user_datain_4    => user_datain_4,    --                  .export
			user_datain_5    => user_datain_5,    --                  .export
			user_datain_6    => user_datain_6,    --                  .export
			user_datain_7    => user_datain_7,    --                  .export
			user_datain_8    => user_datain_8,    --                  .export
			user_datain_9    => user_datain_9,    --                  .export
			user_datain_10   => user_datain_10,   --                  .export
			user_datain_11   => user_datain_11,   --                  .export
			user_datain_12   => user_datain_12,   --                  .export
			user_datain_13   => user_datain_13,   --                  .export
			user_datain_14   => user_datain_14,   --                  .export
			user_datain_15   => user_datain_15    --                  .export
		);

end architecture rtl; -- of slave_template
