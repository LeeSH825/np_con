`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sOz2XXzce/R2EaYLr4G0YJ5hgqA/hvi2fhL3SqH4fGlO1Dfn3vU6SJip2/y13COv
DX0Nh9JRVYJM01QD4DiZn5/tFqUAtmXJeMm4W27WMO3PKDF/060Km1vlG2XtMEn2
5tlO7RjQ7u2nu//rRYdc87Wu8T0YcKCeQ6VvPR+P5C0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7104)
uIqfL1NkW/WJAhIzLc+J9qMa0Iq/f27tdEqourT0NLN1LW0OxeQ+hpNksw6lpEKn
UHWAcNn+8pJniUloGF84od4yQMhj6G7/M+ivs+T9FHlu2BPbcVlgKUFLkN5RMlpJ
VCN2044SBTTrrKg4mIAaCGzvVuAJFAJfCaQgdw+pcMN+JTrWao5rOnvX45+jSgzo
5Cmji7+XMl7hXrrhjx3zsF06ZDz2VbaCbjTDSuGs/7tzHXltqxRO/W3I+y6GxTdO
RGrdmztqHiF8QaGpW3ENyvXf1O7uyzMKdiugxWEbjsqG+5e2yZfcZzjRqPFl+q/T
xmCXkDBpaLWx2yS+Q4fwWk1GlgnRgyp8serYjiD3x8RjtRW5O+SWR1+mzwgugQ5Y
jsPm/jvqYlEFh9M8g+ZBNGaZKyeMYCr3r8tg2p3xC666tiMV/HaeLBEd8Mz99ycq
Czga+Sg/WhaodACxo5W2ThmT18ma82DBOmzHk9Gtb0a5O7vw9qMRTke4kNFhwH3V
YvmLRKqXUJqs6I3bdrbuQrhMvd7Dtdp7ggDkK1Iev9Gay5auECs1XnoWiysnxgsp
rXJSmuO7QEF4/5D/EfH+0sPlnDleBFfh1bfGcTwds0eL057meBum/hO6mlYplXmY
Dg448DLYrP2ZRVIYWK5DjzBZ03aKkhI0m0rod11GZ9SL16qD5ifmV4HHpSS2SLyU
emi9AP9pS3aC1TcMn8fKshPvU+csgPSOVsQ6fNQ+Xrn6FCJHqSspHrj/3TN/MY1Y
Og49f03SDlFqA5VpXFNPUl0Dy3kabCFLXHb4VeAbKGJw9u3lCJzb3mqzKkAObOQu
7AM54x/bbji+gYI6tq0shUPFo382FU4BtdJ9+xB8K+qXuNwWP0sIaF45EPiPdHRg
+6hZ3X4t9w23FJkwY6M8LtLJtC/DHoZSVzYQcnZFbHPzDF6YUoqijPMhgWFFXtTG
EayRJxgO9XrRXBjx10hJ1XxLXdZh+Q2hpQsrcH5XrLt3Kb7yMj4LOMiZezwxCe8c
CBTNp4eaVyMjpiF9fSR/pr2WGh//ihoRr/oyQ/4joEjdvWsgGa1scGyvp+Veq7EA
R8oT8weSaqr/t2f9WiChonHWyt8xSQA5AwStQLgYZ185S7DoNNAzqqy0XBVNLrPU
wkKDOi0pS//x+nrciA3NhttZ5GtJYyz4r4soapc2UKSLkleClMwLre2NWM+66tlU
Sl9+iFFCJRLBtdZrKZ2gROwD1SaLDtHsbrTZcg3bOpxgVl9ZirkOi/FPbc+ziBHN
RqfEo1kByAAsY0OIgwRh5fcpUPU0qlSt3R3R+kVvbMQWEYUB7XJpuEuqhlE10B1I
FHHK8kGYvJQnL5UCpqMJ+P9OLKdJgnosRw/2QdLbTerb0Wo0QsOt/3REBIpysvqT
tqDV2EppFSDJZsV950sJX3y2TGI9hlxLy/oS+Vmhx7eC05IQH3Ls4Cyern9QCehz
B4/fD04VYPkyEal0pkadJzy0lAZip7UduSArJ9AOPsO90bcySV6KUYwIy9VxzSKn
oM6c3WZiKPmdcbEkp+vhxs1A/HMI9cQd8W8dtvTF20tdxmndL2pRcW7qUbYYGA0F
6qIzv7N4ZkXazpIVXQIE4hSDvxXGo92yPXYCjhAGHDsjSk5ZCnBsOduRQe8NviEy
9u2EG2fsGZBPFgXymyysgQjQDAULCs9x5AOwxHc8xDEDB5vGSy5pHM9iMfAFKG1V
JBmJblGuySwZOA/2zBkkHl1KxBDZeoEdjN9ijzOgF36Xin7I//vvLJ8cKzqGak2D
5cEguIPZzp4TtMykerzL+PvGa6GnKWiJrEnwAZH2YHoyaVngzHt5LniCX8f3IXMn
vgQyuropimdNWevbr+VhKM1n89Y/7BnoO5MRE+Tm3FVF+xw66R1P6HdKOq4YPNoz
8wicZ+jP1hz3b4EXXTv5OZJ1Rn3Mg4pfzQAgkIjzPDNlGtjkE9rrtU2KpLhkRUr8
t3m9hnGwcCRAmXDgD5o53PGtYfSjumcEtMNSEfkfzN/7yqKxxhuFolhlXyv2HQCB
nAaB45S0XY3F/GZAxA4QiMPro/qxiG3DxgiTw8vuf5GNeeAgiQJlOBxleMoviLDe
WMkuHGCZnpBfHRMyyem2AYSBiuAsdTDh1c/EWQkWwffqpIh90d3zDQcCzFqdYRlH
UM5aCQ56GaCz9ILCpXEDQyzdXIRPnKWAKJHfmU63ShNXUETIH3pK68JN8dU8owSf
t6Q7aIj4aEjzNfaGsYKUkOoFKKK6RKDvekVTDeFCerWUc+5f7pLogdZGNdMKkXX5
U8Ta29xHx48PE3c5f4ZAA2OZw6cByL9LbVTDj+Y1O/kxqbc9pDbLFEWLfUHZ2h1s
tNbFZ4jbY20D9JrbWFL1bqabNzOhmFi1f+mqjVo9rG/q+hXzNyc/0+Wog2+a0vUJ
C8kvT7dMzXPWvQ/htfZpYCAGZ/c4ewJMX6KaC0mOyjkm8QPWWJz+qskGR+tA64wv
p346rJ5TOddrFPqVoPs/iNdns8vT232OcvD8ZK+53UB+pIQ4W8IU/1II2uML76dP
Ob2cvuPYzXlkMz/wuYem43xGUEqFlI26TXyoo7P+9zpYif73FpaV7ecaQ4/KXf6T
PeRuQxVZs3xXKW/RtEFxfw6NMNp2XfFxWslllbzx7bSY2OkiTXljm+HMHp29b0hr
EGPHZ2MgOkRNhTkhBkZnshTtqFyC/bp0BEIwWGzzrNUkMwLzWXUloJk+k2wQ3LxG
720bH0Ucu8OFUhA46Npw6POlu2+iJNUbvCJL3YTBTKykBlXU7BLfj/jpCQqERSmK
lnGc0NO0U8KheggmMrz/s8nmSM5Bf5d71WRXSqe+MBTzpo2FfBcdKNyjTAPiOpAC
C74DWakaAwheFeef+LC8NVqueQD+yUQtuI6veyuU3BP0/CoVE1Xf7QvMu6LTCKfv
UN7UT/LQBRs7bZ2ZiJd7iYUY0w1CN0DDnzMHgkYdkfjAfBd5bl4gyyelCVKc/J2g
vZZTWnts6uNOqKp6I/BQ1DJjW11LOO03ydCSqUnfaxafsbp3hoVsAWd/URS7Xp0F
Q9QsAdAxrYf6u2xEGRyOfaIBUPnFxWdMOEDWvRi2rCiklAmME6m7G50GAh5baYMa
jZML4yhMxMw3M/0ud4esqurlv7lD7NolkqQQ/wc/urhUM255wub+XAdlS6rBvNRV
B2wLFeOHfi6oSTBepoQkFrPF4I14yMvBP0sle9rSdWqRyK1LgQnsduDbzyHq9SsG
1hsVq4IBKnMr2NxaWXwOnlcUqHKOonIPEV6Kf7fR2ahBIkI8d2+k6vhPlObwvSkO
QbslnZmKmsj4nVOJa1TuvYtSWMTAIzUODnClzXblv99vtLwKpOUGNbKp2EaC8O28
hDrPndvZ3SN0o8hrp69TXu2dYJuvnRghvx9N5PpCKGa0SIuvRsPJ0xDRk/F04txT
oIqNhS/BMMZbjnTfDwe73UX93VFwY85qUSG+izn6LxTF8ZzuRJhbXpTfh6HZNSqD
0gnZgBiIWit7X30lraUP03jLRUVeLcS7sSka49hQ8sCyNpKRGIzDMGsPWZPl0Tu6
ZppktbYclHBLuDBBndXKcZz2U1Nk9xosEJ/41S9wgnA/CFwswCL2zB9WsPSkbM66
oJMw2t8HztAXzEtA8hY/k0bHADxviLrq7KqPCUpsJo/loLp1vkuVqwwrxz3Hm9QR
38ZHwo37pMLzE6GhlZRSKN69x2z07jw+M+NJwqyGV8IBT2fROxnz4PEuqJFUO/LY
wut3Mw3DnJyTezw7zGCTJuaUHnbMUZ3iBVr30rMxYajfmMqx73XWUDvJ6rCwkjrE
jlOUoWrobnvXo07Uhd9jNeUDp4oWCwnZHaVxbmeOtwuWqWR4Kl2I7jFUbdmq8I2c
+FxAX+grwjs9bAQSaPQjtj+TqYNgGFnAqRqWPMnoVQvZ90Oas7nS5+faN3Tw3FRW
5XkExAMqhkFuvtbjYddifE8iG5XJ+PTaHWtXJgT5gZTsjsocWXLEr9FU+AglUoDK
1MFueNiFWWM9bPY1A9zdbwgZglZFqEh1FCj3Q4NzxiUijbnGFdcGMbuLBdiPUhhE
Wy9giUA/NOq8rhW9LAXmSCfDeG9JpfnevYSs05FOKuWD1B1/8WPAyU7ugVuVogQq
aMJbsXDBVHKlQBx8M730xSA11QO/pm0k0IVgLPJGZQlhw8cl9Wf3krwjIeAX4XvN
7ELjpKC7BGPc5etd5kRMYTSPmEvONdT2cKJQ8xOW+Qlyd1IxpIF/lPy6Qs0vGMcX
RirgUySePy1WiAN53FKFoUBmsgU0EGJqD2sEou5ZMvM365eLZYgOyUoWcG0h/MQ0
Qa/SztQAR3wqp/BXycJqcHbEdbW53V6Q10XyH/lGlbRtkuvM2E1++isG/ZXjn2AI
O8lp5EGrTxRrzjzqIA0GGllk3MD18O1TkZqBgKdtONwrIa09wGMalchV0Ek8Tpvv
nVZ9VzLpzEEckyMxyBkO44wJP5J9alxUCFSfu5zQ8tZ30g+VTz+QpskhKxcRIlVp
140fkF7P73dS83eQx5ZlUmM7lr3W6S+jXmxhdPwlDRKvNayDWlntNAoE8yuEUsvR
wViqO+P2f384GI8iKoRXYerYpDP90X4/5yFLTuSJ1ya0vxc7RuVjbpVm6Uel12yK
NwFfFHCwmMbnkMpE6q2K0joppnsG1JO4foVJElrJQLS50illMwl55LTiUoQmuUgN
EPgdOhuu+5H9uiA14c/O2PWus8L2EPz9ptRyU9xBvMbxHCj7JrTfQLG9ks5Sy7hC
XFxB+v/+PG7rnxWD8NPbD/5sewFf1Lb6cXdcTlNbCC3nFsN6MoWYaN2DmnheJ9un
xALjopkWza00qfNFvIPESGXjnHCwMUr0eFhS22RltlJ+uPkTWSEoAuqRLKZggTdg
SIf39q9yrzPzHcIuIoVpooYWmm7g7MwsISR0AqyrNZqtC9BU2qSm6ruYUUx3BKf9
UQItU+cRytK/hM2WGjb+tZzbWBEdCRV8VUEmfFrJ0l3cL2qrxnQeffv8KVIAS3nN
UzAmkEMTFAqCxC+bCKism6XjMtVJhxlJqvFv5NHjSlUS6IKdfxzXdUaXILBWz1vi
6TZ8C6rInqc7S0qEFNk1mnnQQd1hPX+f1mwTMRmEv0HEQpUx4eUgKgTfNJ1qjoOC
JRd3dVlQ0z6PyDmY6VpmBD+vVJlASF5YalccWjD/T5SDzlXCD8jsee1/1vpxw/p5
4KcKD5CUYXJ1y6TKN02qOOGSPZokQGz1bUhAeN+rjWGMF6ZkSb9AVZstsOdmWH0y
DzxEax7RxodExbdokxvnfJIR3HF3BujwRZdDBoH2Gp2x8cU+Bwc7kTzs8odgneXX
5rMM5KsMGjHJgS4kgnwkmZKNCb0ch508/45E37uWpTZwxH07iXIpyKz8mbqPu+6/
sMMdAnovFkxDxaQ2YgYKnnNFizt3YSIS+USP8KBFsgSfjwA73oGn+VCkq1mY65Bn
kQsdsosE0iHdw9r08kliV/lPz6NKS3kAv+qGg0IoFkblxU5CTfQYuN8TSZcSy9gW
RCnMETa/7Q/sUx8nv4j3029U2GUlGi9lalJmeELoERs3QVbKWvvgUu03BeGC/gSh
RKPNWq5hGht9BAbadU9fQiKQuyqoLqvqtWJ74p8SaJauoeuAgbzRYcxIwStuA+2f
Z1jy+2KCv/CLQV8Ko85ix8SYCS2oncgOYaQEXY3BGDBqhQoQcek6Ym3ZukE9L4cs
zRF2JPsremrTeplvxGIGUC3rH7vBybyT/xgDlOFmlLEs85YLJCtSULctk1h+aY9q
2GGAUdCH4L+OruTv+ZmPih1KofquQ8TdIUdP4/QnceFhsXFlL4TIFHiVVlOTWE4b
xRXkxmCkDF75Y3T6VSuZp5KaqWQyzAeU3nL766DALmJvXXyDMjDx/UZHnpQNMZG2
ryB9B8sZ6+ps9KLdzSzvLj7JMSWi1ma8q3JxG/zEGBrotML59vmT/DNRPSu0xDY5
fs6wCGvp+HjBo8M62wD5kNVESGBeX2/YX7GfWkS8ekuTUnqHLSO+hkaU7IpcE5mS
DeP5NmwMzupKglIz+zY+q/TFr9F6vfEIO2pHYKGPyAq3xZUcC0+X6TU1Kyx0Y77V
QlxnOiNXOI0/O7BMcteBm6avnjPmYxPTupgueVND7Aqi8R5Fm6ZzqNU/j1jmnuqq
gqEULw5Z6iqazJZ0ycRD01nMFZCSmFrkmkq4j7oJAagNOBVAV3qTm+PZBIw2Ln7g
Rn6vJvqcvIWvKbA3puCp8y+YII+825G+KF0eaLC/amg/aHcqJ1vf/BHNe1vQf+sr
dPLhCLYFgT5bPfEZ15+f49sgOM4BUUS41LukoNRm+LEZ1VtxDGnIA3C9xuk8Ee0G
dIgU7Z9W7FKfDbFAVx9orvd7FV1CmT0nCR7trBhc6eKM1JjnjRjXvvTgbVDTodKu
1yGHoq2liRSL11oYFErR/R+y39kEjxjOM5a9fdFEH/OwT19MuIT1qfweQHH72ZNk
XZSxWZL7jf9DW2O67jZ0+DvO+e6/zPkxNTs1t2F+nX9jlyFdNliNNWKyvD/XkWI+
hEm69oSPrM79J69gvUzv1Jle+0nT4gQyRK7Y3K5aHTp6ZAnT0IzJFakiWDUUITWd
3Z7Y8Gfj+xH0f7jgk9z6yx0zxzUbk0ZxCpUDMTxo/RTaj9fxeqCP2ffQk38K8DQa
IjcuEoFzXZvu52bCMumLFtzVaibFEBm35yye+bPrTYOlZY3mJIGlnAwzxFSo5HEa
M4wmuGiamGJsnCyKMMajtZQHQ2OkVCpQ+uCdiUra6Bon7ryiv051eQUmmsXoaLoI
gpaf7KnoYGYJr1GVImZXgpgfDuMWYNw03PRZwFxksyqWS2iMoDCzQbkW+niy26Ra
hf6YZGPt1fzamwzaF5+iqei2LUTYy13rb5H545i+GFURqiTu5vZ2J1EIgaF5Qgz+
im3zSIJKXApf0hQgwfzrTkAP6CezgyEd0VRoC2i2PG/WJGGAgYtR55vgP/acUmu3
w5p0COMCdtxjmzaVUnKjj7kTD+KsfafcdS0sMAAHkL+K5MIhkbMeILOh2AwJijn5
hnU8JR6ls/NEJDAdf68gWFduehXAUIyd2c5Cuy+TGKGqR4of2iwzdLs9rclPpNUd
kjijbsnPQwbh+Q5JKhTyGzvnBllmpxHKrSNn85apydFPn0gRt9qNc6VOxw1l8nMd
42REMKbIW5yqd01wCniY8XOV9FcADpm2umwNucrtvuCqONBE3uAJnP+P2eLcdS8C
uzEACrY2YLFBs6cluCHQADZMCIeytb4eiWmLRavPIHndFr3QiGeR8MyQJehWOsY8
A+llNBJJ9aNr35+3dq+7F7VeyyhioccQJEf8oFSEPFFrvF1alreSl8KvpjDFVhwW
hJPE+ZM4b57jyz+1JUsfnekI77oEUCvIPkdcPJpqsZoj+EqAQ6uKFweHteUxEjgH
45UMzTpTsp7gL887w3cfc8RHbRouxgL9X30drqC3NsB8JAuaBQ48YcVvgJ6LesNZ
RJYuiVAkCgUGptFxCr7ucAPD3pXVhRNjxdBStKQUjd9OsO9hoLpmC/MLqijGyinV
fv+yxtWlWhxcHpD9pIe6KAscT0bNhvftrxW5hU/M2gfJS3tUUMAhaXPTTMFxaw0g
bmICXbqErd4xOku84i8MaoJPFMyaw6rkUUJmXAzlplcJ/b2SAdnKNpbrS1i8CAqr
9Hw9cONDjvQ2dInuSUnPiI+ZeJPlKEnxKW3AOHEk9uPlRP2wuCM9JN8AG3qJ2a9G
3C0itu6XphkiixbjP2VLGsAlz7l2TwdoGYh3KzoC6+HqSa5HEmbCFVBZQgsAtNiA
IfpvgPkujU7xDOQCFJZd6AhiOY8Em9MNHSdgGQQdG4idh0bVmUgGwPzT2hbNhamZ
6Qg3hvM7wYy5aComa0zj5FntqeIL18rD1k270PPCYHaxcLbkTS22Uij0Jr0gtY2V
jlGkhpMbFnyaEfVVLhrEQI7IFmK2+8xSj9VWDsbb33/z4ThYVrFsoSUH3Bc4bqK+
4E5jfDCKkOE1ic8YV+kpAbO7I7RiNWFkPygWIKpUs4RFC/2WTg4xcqdx7LOKkMFD
s9n9NhIyZXpcY3YPYI1+N+8rYVKH5rfKQQ06oqS2tbkeHkghW8ZAx9lQ6SnONDrQ
3hEyaGY53igHj2Q/klgSw9NiuJ3+64GBtVVnzRmY36am6klFptPOk+Msu6jlEUjP
VP63R0XRlf7lzRY1vk5h4idlNOnQqWy/8/B9vlFe5ClGRx8ZazNh+1vM24tyYad7
QI3xdaO+r5aN9sToMj7ooQszDzqmC1d/rwT//hnwS4fU2ht0UCRV4GG1yX9swHHv
ZZ/ztbgBThb5mK02NiR7uaQtQXRAKlEooMyYTmf8vcHjry4kiWW5bgQjQ2zL2j8u
naY45kgBU5aTjwPXpci82lBnv/Iuto9bke7kzB7ookAz2DkAm9K6AcTs+Dz1KwjH
PwaPpkp5jURogu6tUgE+Ov5ZGfK+jysrDgGjVbF2mUdMFVW2UgwTHsCnXdTXF5ws
qD29oHkPkZtk4sK1I45pdezGveH0LojHXNa3ECf+qmo3KhilzmcqKicIPjEpBb1c
G/uCKvYNyNCiUsH/t+4x2upbn8BM65X3s6RAU/7ea+RZU7Ez1uTHNjVYzpC/PeEo
xEBB7ZpOgxjVM8FjFMJ31j++TKhTg/ufn/L2BRW55H24j6zjfcpHu2axwH6/eVxH
AXolbZ6Umd5HDwrdtLDzeSqpgyCrBxP21QTFXjvXFvgmEDAmvZn999SbQd8OAZFp
uKG2fLlTQeiVTtzWF2tl7YPaBGjgXr7lYuyUTsfCDXXOdFv41wqe3R/QLqG3cjc+
xPCAo48lqYoyFlkOrw7eT7lrqAUWSkdFqAi83zlf0cvjq6zDlqyI2a1fxVrRx15r
dthxWSF6+Cy8SFGMGHt1da1eff3B0iplyWiL2IXhID1jRznkW1sKDObZcGqYxcSm
1x0CDQWT5ODr14SD7xUA8Y6u6o3tV2MihIHUegBtVEjSSUgy/pz0yJQ3KVZuYhzE
e5q7RlXo382s8AfqHeK/Yq8NsvMiWqxaIdO68TXIFR/jLwEnjOIrYEXiUkol5L1T
fqQzoVmdl2vFoQXTpaBN8Nj2XCcKPRCUkpSKN5e9TTdFxN9m2sH/5oFT7wXd+Xck
riQEeb/E4G4QAaOQE7i9ZySYJtW3JSdtm2s3d9XoI6iiQuUH2DIXNpNZ4403Ocvh
qsQ/pIY8FrEkqCgodlQHaTLB18KOdd/FiBU+Js4nOf0GMIRRzlE8Y/6juTGXSSOF
EDdpPqugQxK1zuCKeKe0cH6j+YXq6L9U13+r5FaGDueVkKrgUfjEq9jejwWcFXpr
a8ZyWG8MukiRXUvPbfx1GQNmxi+eU2Tz09HRV1vvlpzVjq09FuRGXfeLA10XMg2f
`pragma protect end_protected
