`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Zwqu9ukK7UlIFDKnG1rr0KLHtl24Zx8tsUxFXHMGyFgmQW8aKd7d1WHthALlq1gF
k+aYTcvWSABb5YLdjFx1HBht9vubkddOZK8W6Clycjn+GGJSvxi5JjKEpPRkD8su
DjqWG20qOUmv2Kf87PfQAtkar7lw4X0olRJy620h164=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21696)
Ep1UnoVME0O9SWhH1TArss/ZjRDhU3IH7yOdGgnLebmThlEWegpeY+4FAjsFJt0Y
D5KKcc2Hkrg3MCyl+gTh/MJmy+fnW94glkEjva/QO5E9cpdexiGH6eosP1ybhTNW
WrJzXMfEa/mdEELTzQCS9ku6KDnmiINs4zWtulx53o6OgQQ7Ivzz7dzhEJHtQVyZ
GcE8JA/0Fgn2XSI0H/u2H0AfPDJ/hmeTJkD7Mw8lZdq14X0z0oqDywTTQx0ECJKj
gbKXqnz2nmSgLpNHHdcY63C8U9laUr96XQk6ID2cC6niieH6BBbrh6g0zZeQFI0F
ETIzeWinIL84krImomRwWopaO1m/s63LIbBqHG1muL/j9YTJh8wnTVwIUHRv7znz
hRpqMWBUkUZ1ffqiGN862pZIJOlffwsA0+xjkjWK60lP2mI3y2iSlf0s+zm9Zx7O
4VRpR1azUGPfHjYJkOuju9jx/TvGeVK0l0DGZLogGH3e9D4JvX/zy1kAGvPttOOL
iK2OExxqQo/AbVHEjinJ2SPQyNMXoo1r1TNNlD3/q3nRu1/aT/1GcsvHQD1LmFRu
8v5woVd5qdvWCfBnKSaveBCo+iut21yITxJ+SxkEGMhT0K98FiuV5RNHoXjIUKz9
JJEVSH7nHxXeA5I1qIK/jnW4aBEfeZ1PQTuqi4HIGJ+f3Zi0TlF3J/k/EYjhEw6K
L+/O1val6iepBcgI/FQUPZ871UMYBrQyeVJQbM5zJZlObTvpVQ4MU6m12k8X9sjj
jiB9mba2yni931Lir3Ikfvj7sGlOVwnzEoI8zxI22Lxq1leitoWg92E8VJDHbF2J
LI4eX9H0+Yc2p9wLFtO3NPqZ0na2J4yGfF3HYmnfhWFO3T6+o3FNCHvRD119rcIX
7E8hRrx5Qz/pak4wdDXaloP5/EgBUyFX7KizkXZRfLZ7SheEpHiIA715j7CjoWBF
7Kep7xUMx1W5Yk6cOgNTTxSVuOYLsc+JnzFBjvhy2Yn/Amsq2CHN2O4kbcq3ETBT
vwib3lqRmBPEltJwhw8i2J8p7g3dJ2L8u/d42BXdf7kluFcm5kly0i38jmK/l+Lg
8ruzt3aRHPmwAsEQaPITTnKEMxT/DG6GbfGTjpESRljWdmzbmxDp61ksHqwDTwnh
ZLy0ZqJo/UnKySrphO8sLJqsnTailpG0Z+WJRoe4nblEeyzaLK7geh78XbYMPtZI
4LT0GX6xw65TEZiT7434rtuAy4QlhmebJd9pECSCmPEMXPJlzMBEMViXQP2Z9NVa
uJbgTd+B/TmYh/1LnsgobPLGK3TaNP7lEwK4HamKePsa9W0By0yYJLKE1u0KiyiX
jnxBQy08LFfO2GqkBeXVy06AUVy3pzY80Yy3YZARbypYpUq5ay1+wxOZkUAsderM
6ShG4fME3mG2wptR6KS+MDPQgWXD4HazjvPYPc1c/3E+1lApVZMMpDA1FDsgReTn
Go+feJH1cOfFvkcxhn8UikXrnoAKtm8EDp9Vl//y4AEDxJJvLqv7pHLMsPpFJ5aH
zyVJszZEyb552AzKHrExYH9pMYv5ENANgvwCIsNHEtJ9Qw3qihYlu8isJkxyzM91
IF5a/lOhfsWc35LKxcB5LCadYdbzfYqVv/EtL0HthnV3UJELvviv2snLbMv6490t
zPthh65zwaQJP5TrLdeJOw6buPEWJwZUKtNObQYOFGbxOZ0e77xRMmcl/YM4lVFu
6xwu/KZvSQOz4NMiIHOxpfWmSK+LyLr1kentkHrv3oT1vEAYa+s40ZgNcUQNTvqm
VFVj3P6cfFBcpCwvk4cSQqzIHQQAHYWFz0BpWHa8yv4ti8WWhkqM8Y5LFX9FpdUY
AnNRPm793fDeWENtXjslzm5jhnBmRoCp/wDC9b7FkPsOJGX3NcckmDg6opUwHTyP
ThGs278LtOC1pg5VJ4E0OGdz9Blnc0kKiuEwcQo2zKSiNLLMixkb/qwzkutOtXGW
GmcYxHktVMdfZALK8veyGbRzXf2VnDFpuJSDmAx9HgXDfijMh/raFa+fNPH+A8QS
WmsSGcsU2uuFx3zMt0JtMjCXN4fvxtxbVG8CRPvQiQXxN4WK1MTKqydhtTVszqSO
0pO1BNc3d0cFkPYulAYf1QifkgnWp1KDkNhnyGnEiD/mPUr5FaZrvE247to9EJ1U
dumsbu9ALp73HRm0Mhjon08SqBL17FPLjzYzZk9ctVy0BkI9DXdZ2imXqb5HfpWS
c0NtgDpTy58Bla7AqE35cH0Al11EX2DwzyDauDCmP1p+dr9UrGOE1YtFw4NiAbIV
P0TOwR6Cm5iB5txsr8KUvgu8wsHo2XIBSsdA7OqS30koAsu+LN8GgnldbBprug/o
XOjX/j7jMQv4ttf5xohfXI4+4775v+3G0Au5Z93ypbOQNag8pD3i9xZ9+T0J1bO8
WJhjjmld4R8WnS7OA2T5LfGIOMK8YdE9fAbvRnWmJVEBgxRNrvOcKJWW4lIJar6p
TzyYQI8kJvah8SHn0LgUUnjKRQfDt9gIYscxISgkhCTE+zr7BalfCsQuK1lZHkc+
i53D3jC2OFwdk58+yTwPcj0YcxH9O0Rkz4JCfk+mMErtXXabI7nIzFF5T9sqyiPa
gnMOGXd/WOhNTOk8aE3c7h8y5NOup0dSE39mcdlFD59NtAoYUuckaPcFQs4k1IwD
uLXq8gHXcC6v7sMKgjRvIMbx7ooJ/wsaOBuaKe35u0houIQ+2dJRnTbYYV18cOUc
UHS08lrXBCaaE04woy0GBksoXAyw4B4MQZ1kNNVwI2QLykQtqg2wvnizjc8R1nLT
GTbkqZAMwelmr6eZDYjXZ0eTBL8ft9jx1MvRRBTjYxeQ1bSLMjOKeaYOHqtoAHrB
7OdkvG1Wtm5pnSr3R9PwX+olryoRYpbSyEpuNlkQcOAR3MGxgESHh71+JlAH/09F
pVcMlB7HJkl5mkDokWGBvXwZomF7fpPEi3FWhdLGRDbaP+3zJ/HHqZoXUp1LtX2N
gBHjJKkqPxGCJU5VjWRQZJ5nONX1IBctIC3Tt6Hy8xv78q1sMUAGM6ECs1RZ3Drw
YboIvA8HkLJ48ex1NRjkS/Le8Qas3wQyrOX2fUUgN92mRS/UoyDja795L3chGJIZ
0j1mQ2qUuF/TGz7TiIUrNw3HDy+By9MVtVntFrkqQRTeo9f9VklPPVZlvui38Pti
IjaBWL097Ivx0WWzh3Ky751/sQlsyQif9DzmDsyVDEhSTzWpj4a2l0/yfu03XL01
fLcuzv3iNPn5oPqCr1ckcAF8RvTvHzhyvRQT28XkcikATan5nG1dJ2Xrsbgth5GW
WRWtXNpJP6yQQ+n54eLWhv3Fm3kcjVXyRTumeC819P+j2mN+YQbuxhsZUNScKplY
RV0n/Q+dE/b521KeQoHlJHqunVYSMK8Muj/c6g4UXYNqA/uJBX7BFM+6bGmNEW0X
RbK+8h4VxEoKutIJ0paZhI8dI8nlFIXf6UHfTq+NWc8fRmXr2t+UWUhA9wjtVhXZ
ToZsfj6MJn2i3n1bEQroLtWXIZZXW3dgyJtFAbrJCeJYguam+cuutq8uqs7lP7gZ
xBi1lVJ/yYr4BMqQNQvF7wMUNTEVHo5qM0pIAlMRIT2zH1/u6RP+42SVocO1sPUI
9RwBBftb/fOkCe2ESjT74G5i1LLJ/wf43/t3CsaYeYjQfwCAzuZ2dbpqLEf5pFGW
bwCHdyca6p2yWqdlA9Kn5vXJYbXnrIVYPr8Hl/cVQ4VHGtJLG/+EiD6SesuuYXjA
FP3LM2vhgD0EFmaq9ZPeJBlQBly/vInvhz135dHxUMcL1DNYy/XdiYIH4UWBURJp
TcAEOpj/RuEp4FF2vAKJo/QD/QAqbissG3zNnKStdxGie9yK1l0ah8tXV/pBlxsi
y9EOgp/5hgUc/U7Z6ic+T5sFlHh4tp69ICjIcACIs3sTpaR26YKZElJGcfbIyjJV
HUcFxw8c69Vrf4cQ1R2/0pRryElAdgl989FuMWZW4JZl5GTz9eoT/UV9GEDbuBaR
mdnNigjQLOsYd23CntDGMf1sPAduaX0Yr6FaQRPvOcfG0l63ja6cPDk6NYHFGbry
4Js0uRbTwBVVQWte0+7h38qjVNTa59D+zodkhLia0qEVzncnzpHuRmFAgOXDGZg1
I0hxj+7AFtENxnsREgOdGaxURZ8mhsgkkhYPq0bbutbqouZk+b2plTKqICRB46jg
asEEUS4sjXvLT4UKjaO+sVaMAMVEVZs07XGcvM3a8q8bdnQlR0nEOJsPC4iZV4ri
1rjJAIveKol5D6u03BLuaNV/6X7TemaXYq6wn4QvPKwoHn2gm85AB14eKoWrcHZl
pEd9bEK7ULxE9BgZhHO67upR6fnLdOnjJIUMEfbxbk/jsx1wc+v6dM7FATyj68fX
DemoO/98JyeA6gUo/wcf/0BB0cY/dvk+b3+pEYAGrVtmnmN0q9bKuAlfhqovaiTr
CjNy85IGZqCdjtv4zncEQFRpCE0F+oAU7vekJYGPMzAnGIufHA2MfHw1BgGQVrpM
st2VmqY9OCeS0+h0PtPVDcb+k8ZMliK9xIgr/Z+YnehHfpre+pLz/WjGF0QHpwo9
cHhuhclEseDh8D2mZJDsAKRRCs/eANErNr4V8FPbs/HS/I7mECcIue8IbEUtK4Qd
/r6FuuF8CuIbZBHn76Ap9Oc9zanX2VSaGyxf12NeiRjguL+8rLF9uzRF07i6Yhek
y+aQt+JYwIbpfWTlzpxonvvY/ZS5wOuXo7OmI0NIZtiLf7D07T2RP4e+XrdjrSNV
JV2pUMjXFPIENgf+WwUQIMoZdgAnVEMiXNiyS1lffMzImOLCkgGoMP0QwwJX7/WO
COgVmArFFfJl5Wz8iNVXhpv0+v7qZGbeiJ1ZUFe1Tb4nI8njfYiytR8Wtx0tyIt+
CXHdH6Sii0LTw0nIkx2vrrAF4Nzne9eeoDyRMzmE/7zPN0FDApxilPfm45fJc++g
lbkA7hwXJ5uiH64nMgsfB17QP7ySDeivOTa9Hx5Z3ddbO7JzOAVEqXMFrNufYyNJ
NnQujNS4228Xjx32aEbfeCoSnclzK6dc+ktCc64RuzA83joA95Q+cGSKsrnD66oU
NU1fv38nXVi6VqsRF5+HYnIjeBpt43K/bWIHdT4+rTcSCXMGGUDn8Ncf0f8wKjXI
vcHI/xqn6JmriTWdK8i1TXcEH6N36N4ns6YO8HDMEZvBI8SYhVzfPbD5ZCo/MCGr
hXzSV3q1rG3jVuDTFHeOYGZTn2mJZ2D6ulo/XmlUtwTYtzZbEZtUL1Wxve/U+SRL
1R/AmhyZ5iVSy9NJP/3e3pYm9gf4I9DKUXHbeFjcU6BQW/cvm3D/fAqJ2KNVj02v
/r73PcZ3dNjqV+F91CxXp5oEG5JKNkdvVcpM896xwqqOnf2CNon5Qzo33i//wqdE
K4sa7+3862FtjnUsXboITXRyaYizw94BGR2m3T6UAwEJ3KaFziqRzqY/cXgYf1+o
GsGa+QEBrFNrtHxYCWuClOUQ9X5/ijud9ocCJ+NuVBiBv/QB+Nhz6mYaoG2n0MEX
gFJ1jI2Jx8paZs1JXfD685B9+MvOOPbS9q8ritKOYwIlEk5DGZFAz/LvLLBkUyR1
BY90/ghwtwvdPtU5NR00dDvKhV9Recxry6j83S7lYCfwpnKDtjlBEee64Y8jFVgd
GowyilyxtEI0AJMIOP0DR1VNgyKpWoCgDXSZJx2EyQBgFhg3k0YRRslxA+7xf+dT
ECQjpHDfaazoqoTg67SqEAK/gB6pbxHzqAFY5L0MJmaw8FcUjD+a5Uq3YSaJ6VV9
5HQEVx6aWACUmNcK64dMiqYToet2YYZnAO6n8sC1qMpCThe8C49KbziWyewimeA6
av07/s3Re8AWs+ZmVn7Mqwv+qFlGkUfs7HILBNHp45Zlr2NklLcaJTMgdJZCufDH
h0IGxrhMun49om0a6C4d5Yr5fx+7V+9SGwjLVhoPgDvjWJJ0VOee2RgcONeWWO7j
0vaNZ1JfB44gbxXlI5TUC9vvNwEnvyDrbXEa2s89hTEoIYxzIb5SqQqSHnfEJk6j
7c9SzGhPWtviFfdt9NDftzUjFjcBvYSBATaGO6GGnF9qPeaEJX9EJMFCP/78VXAh
kwPnAEJKNQZ9XJqaD09uskwXc9vz2AEHubDxRy9QMHrkhEA6GWt0BpLgeTyZO+r5
g4tNkZ2DQbQvqIoCSaTwb6KZk7ntUROEYMWHeIlWJDFNl424OgcEYd7nOwAieLyc
BkrFDSIAxCyz3hOCDqJlDwudof6IqkQX0Aa5hkg4iDaWgA0mdy0QZcy0jjDWK2yO
7Kz9u3O97OXn2fydjVfhzY8RSauI0IhDMJ428PQEhDwXpD25vyGxuuBbDIw6rfW5
T3hDF0QqSiQHl2rKM1U0wFOXN+tC8DH6rEUdwlbH2MfAtZ/oQW3cw6Cd4G5/Tsj7
Sb1RLA7G4yhFYcvtV7B6nKlsySBumUhztsphC68mdKCUhiJTLxe90xegiNoTlkbs
5ocE+WC2q+aJkKF4jDtTg8G0SpomFktam9Z5s6lJDoxpW6853dnw/6NudiAjBiUr
0G6PqmuQu/DjLRZxdPxqSp8ytbZfzh3VVxeTzz/Nj3kfswlyx3WBrac+tjj66ULw
5rVEw268cRHgzUv4nQ3q3IuxR6BODV7xQGTuCznxyYRPOrdximeXwNbMCdC3X8hW
qie4WXRVGrUBrrpvoybEripZBmhf1Ewfr5Tc9rJn9pHxxpU6jqJTbyC6elg+QRt9
7u1ms2aCaEOUOu9hqzZXqaLbr1CvpXx+C3gg5Tpw74jhHwYZa+TEeeEU/PwTkrpC
LYTykwMi1sIXz6aW9V65uYUyeqE1XpTXUvd1QIvqBgv6KXeaTDUOptM+/jiZIAiS
H2ZG2S2rVY3oU7BG4yfcbd1jUmx2KsA/DkAZPiwr6sZ6k+UW0LyMf6wR95u4YrUW
9hy0hrRAZWoGUGwwP/almdCg9H66GDQH7wTy8UV/YBRgKiEiiBZkN5wuzYacvv4r
sJ2mKuA4hx9fIr9+7j6PunwSMnVdOdlTdx7UnRsyCMt++Im6FPZND1suYX6jeXB+
FPugAWhPw4v7BodLlI2FDC2vTFCApsEbedvrr0y9eMg+a2vk5S9fpEbwB9eP6bGS
67UDO1+PWk8I0tTE219S8Af+4YyG89wLp4RngHs8pu0CV2sHnPWaiAXpWXbJOyyB
g8WEALTumaGK5oONjacKFXdNLId3FBoZL37nKuFUkJP8lE5KQ66hhUxNU5DN/CRZ
oRuWPu5yqHXTmLhi6y2RGQo14g0Dg1iREIJCvLH08oTgw6iz/l2ceyhB8wERwkT2
9qI18gDp3jh7wnZds4d2hZY9tvXRRTMk2RSNRoKEwX6n6EA/w1jUgCPnC3env1AV
xYivERVV4ffTfFOX9QiP47awPTuffaAGNvvxpxxlEexKDzR4Jg3ZvfZ6duRpKyND
5hbvLle6XfkM43qlgogAo0irLIMOoC5JY2CSYFFK6uPyn5GR1wtNP+au/Zg+navI
Tv0RAiwLsKgWKdTsKQL/yHzxeEvIZMN07lfU/aM35W8+5OuZOnf2A/0kFWueEE3i
ebcoH8cmTxfTJRev53lKhoGfwoFTBHy5K6dWQev+ZffbjBsem4KP6XqeXLR4C7pc
MSU8rPaOXglH/UkGah3nSv2hK9YQ3DBeUyfBb0xiSS6wljM9/oo+wa3oGmOtUVCL
9cG22XOeaSgxAaCVGXZHjH6F7uedq4Tj8jzCB8MtSr4LT01YCffXCGLcZwbXmtDo
sFbKIzcaJtzaNICXgjj/izvQ8HwBbbr/JVtf4EFW1G8oSpS8+q8qq5lLa8J8gUCo
4gI4bQNsDndmLwFsML4CGIVaZYrypy8Gt53wKvFspDFuKBhzfpygIGX3flzcjwtl
FJRLHghK7KF83vaRW96T6+LQUfx5l5CM+iS2E8vPTsOo3cJW+6r44F+seFFVvy8g
VmpWNRAxCnIFKdLPWptOnd0dcTbtogbprQ4xCIojvXuvHSaln2M5hRSR6FuBJt6D
8JPhfuMeVdvByC8D2nJNZwZduu4SySeaiIaH8UrOdnzAMiVEzSLJDklx1FxI6zO5
v4p46rreMoFfLO89U6ZHdLvl6O7EEf5jCPhMthkkteD8TNJDxTXfTmKmB/jUzprG
eDPuJIRFdeGeUIbKkVjMbcyCcgpdefAcw86zuq+ngEw8R4jEQ29TdCZHUIDZq8Hj
D8pc0DHBNzt7y9bIR6udBn6EaBHRJux4DT15YnI6TkBfrFUknUHVbi9b3YwxobZ1
nc6HfP/LFywAhowEtn5H+g8c/mdW3mvdukVXpC3cQu42p2RWn5j78qhE72fLfgDo
1OUj1o/Wa3BLO4p3HHSEajdazWzBctk//YcCrhxMb+SbKxc2Y1g/yrFCt876qS6e
nbxo4qoB8JXVo9jrMPj4H9CAPQAUJ+BAihOzfEmQAMdBOiw/39/LasY8/DU7uoDh
HVS9qwcFFko42SGpeqvJwrMZF1Lze+ll2GxUciJulHIpBO995xjxaFoQ45CA6Zvz
C1psl8UAuUkDR+HJ0JBDjoWv9i41ogoewCI1zY4SdiMsBwR/JN/BrWKgLwmMjpYb
iKB7tGcqnbS3/P1WjzPtRwrIkhu1IgmDLY8Fl3gJ6ECqjMiyTRS/LWp7jjdOBgvl
8VhHVMDzDYaJp+cjxfJTdfqobY4kuCMy/4PFH7/JwoRQ4kEzboF/YYphXNbUtpyI
jHrwdSmiDauh03PJm0Ch46ALWGOxE0JNLRbvBq2VKArSF+C/av0CQG7fE0L3SLzj
UpVp4fMNU/W7WtCNK4yWVRU/he0Ic924CoxXwX7yCxgGVhlwlrMobSdd3HtjL+2T
aKcNTpFhTsVbfwS7cnmwDNGt7qtIoXIC9x2KQ+sasMUWwyilRWPhXjWkc9E2hfUK
PbP038Zh0KwCIPiJ1Wc+wucrrc430B0fJa4UdCrvB14C5bu+y93xkbAVGi9gmv8t
UpfdF7BuQTD7hOgzG8CzxcRDnz4O82dgZH2F30NLqXKKSflmtfbL/AHvajkZR+OR
h9CqkR2Iamk1Ja2nkMV0lYqXa/1vHgizYmAkFycO+yu/wBrVdmMans4VS7fge6Vs
3sB4AWsl0uG7X7X11gViEnkV3L3445UmanqiGWB4/lF00Q2fM/wMMoNqHNsvwujt
GxPYsZO4oP6afSGEXC9Jf/hWIsCiThY7LIjrSW+O+HPgDcK8pgrivtOgiq5k+K5H
D2fX5rZgbRWzWjOJqaxeC0hEGDLggDunjm6g5GSXmePXNZ9rUYL5V5tLT0YPPf07
gXoGzn51eaGSGv889potMDfNfM1S4FK6qvbfJDWF4XUOgd+YT7vHbYAesIsowm2X
cGlUXp4l8cYc56+WEeceoqpz3mdcn0/lP9y/WLWiVbyGQVE37rVUTTPoYVUnNfAl
A+K4X5cd9uYSb2sA2a/NOkMzZ8l18NHUNtmeOhPfflm5bLHSWgLLj+14XsPmr8sE
320fH6CGwGXJ5LTvJ2VDL5a3IVhZVUXDP2MiSBmpM69dWm3DtV0U6dcEqc6yHzbr
ywpG24VtJXBSLwcj0K8R+CwqkLpVzk6TmSNY1TVNQZc8wGEMypUzIaF/s5m8l4rE
poPkoNroM0zO61XMlj5LfYBsOMfoz4AiVSfX3nIP/WO0xfQzWhuDveQRjx2Bh3yR
/LHRWWjkZ8xZq/SiIco8MD241zobGeOmhuxGRjuwa200i376Nx48gVaGrtFE02i/
krm1meMB5OC4NnFdPPu8XwktXj/ApIbmkCFX1x9DtSxxI3aodlOmwASEQ9rPgobm
/Dgw2AzfghFrimLpBYU1m95DcidcfTLSpgZfbnLrgn1TdiJwWU6TAOc35XWvs8y+
qBXG+V3/xVrGz2QH5MT79xw8SBr0SjC7+VtC2J/99xccO5zA2B5Pj13kDqaUfd6W
eTxGVUZ7RfhR8m2aLEsVWlrwT92/r4ekEAD2r5pqNf6LYZIJNGA89KF2Hhqe32AO
OY2Brd4vU445FjDP3l2jBjLO3XmD9p6085X4GE1kvyCfV1oxkGnYkjSRh/eW9cnc
RvbPkEABiNFxynMgc1XdfFe3UIBha4XKAk1yz/d0c2CRuCtQBbgHjOs26Mm4PTJa
tVWcWoGz6njbeXRpSfaFrbiGU4nhltwC+NqWk5IwGNFslAY8jo8zLCg7xrW+NoY2
LvWMMNeUn0GuTLZSZZn++AhY2kzJSCZneYTZv+N9jOquHa/DHXwKhaZNexGFJe32
d934Na+C1B8LIQgG1pl28OOASmCb7jLbvBbEZbFbTiXDH02p814E0dFysXeg3g8J
grxIqop9pXAp7m9rphmqmsaNMFqMFv4qB9v7pDcSUEU/62VKspDA1ba2Q7ircG7K
xwR6kYR4dW1WXXrDguRsyZsSH5mF5d7sMZTtUUWUaGaX4GnGRuMlCbj7qoMHaoDO
amtv61EkvVi2pB5w3jOvCoKm0a3Z1VNzGktmvIrLlKZgyZrDGZm8sr/gykldQGj4
QJu8q2/oerxcuTUZSMAlKWifxPLjtFEvlCXozhPK69osWT4iahwyS5ZZbmn09Ec8
DUFZPvbZzU/ezwdpyTc2DpFzeOamFvf/ryHJOozQK40KrHwaI/klL6GtlxQzjwiQ
9+UOH1BxyxMhfNxYNisdwfc1KeirIBw4h9fRWZP/yq2Gy/BciGQeNRyhwfTo8A8B
7/eQLb9o/5D15aqUh6WThVTZPVCTmjuXar+qEukF4yE2CQrlACOQWe8TeTlFjYew
pAJMIrig1ygkZ1zbSGnGHV0OOh7v3ePwoC6q1R877O7MoatV2xDnrWl6EqfqzUb3
T6oqdAk91r8nQc8W/ZVuCMkiZWewFGuStXkxcyCAqaNMRDAMpZL2YFUnTYBHP59K
aQJceRm+l035Lcr9YVsQFng0TYM7BzGPYIpmLhtDhnULSCzoKA4XOTLNYEuWgNcc
bVoa9kjKNJ61kNLfmD78IttfUybxffO4sI0PSpcRerDhOcUfp424GQgwuHXeVIUw
iLd4bOoi8dJGRJVxrvkpcdolA1BVvBZaghU7kXeFRme9c0mwXkxr6Z1s4pu0BEr4
TD2nfYRtNLgxsMfuHuhUx3qjpnULfls6XqJag2LNmWqEax+HpQ9W/APtuJe8Fc5K
JYdsnv+xuRLZfGddIt82/lCKucfX/13KnR7Mga1H4BQbRiBmDd+5khNUHMIN1+I8
lLPU1EpuUIjyt13Ot3r0BFOAMAzxBWUh4Jfwf/oPYE8+kbnd8Sz1WEaVbTbB63t2
AXa1i1H82YuAulKSVlCTtfBf2OpLxhVO09erQJmubHm63gTeeI0q4UqnMn007S8N
RUQISCCeQqW8nKhjYONE8D2r6mv8fYe+C0EV9xBja+e3zKfogkRAess5RNnHe8sm
fNZTEwXOe6PkYriDL209WJKSs+z+qqp59Sy2XLcQ+ydPJccPlLHSgtPCrkJPGahB
NeqHbMg/5nc3W9ZDIOb2YaMy6VpVGneXv3hSle2BLRFpRGz7SA3OXbR6AvbwWh1X
55nJ3SL9qadKFVQWtW5ThCZ9OnKAes57X6F761v/wqVQE34eNm4uLkchMTca4cas
i0N/jbIJNqCF23MS3Sp1WkNbYg/SQAPZ/yzYsm5fPO8o97PTE7MpL2/e9T0SdIWx
qf9aAvC0Zwo5Q3q3VvQsASdp15i/uE+qMn5cSzx83/+2/DvNTHeMNfsgR7UNUhLG
sDDG90euq0NbWFEmFSurBWZRBP/zkczvB6BiI6kOt4aJ8Ts+gO+0WCHhxKUxULPT
ErpvXJRTw74GCbiULzqEsRwY61TWuBPEPD5b1q/alwigEBwWMwhXyB5DO3LcU3aR
nrkyfJ6dC1fFLQtRS0hCZHh2j+5HXXl8M5YIXEP6ThcJ/v7ufjeG+bXaASvXubVB
n5h/HedqqolyJQTVRnEcbN5Yn7Okd6/U69wPXnpahSGWn4vX2O3Znmc57MEKffIE
GhEyCQicQMb9ibZ2ReQUzp7O9WHdmg+ETjXuqq5c3ZI6svfRberUkWIyKkVukKqg
UsZxnPyvZZpXKMlGhmX3Q3V2XTiqeevJV7v6Tx0XhwTciUL28r8GFxUDm+CAYDRY
w0J+viq47+ahHTXGqWvtSs3IddHoceglsN5CG5fozILfqY2K1Nh3nKhb0zIUeWkG
yugrDZGoDx0vu2tU4JqM3DX2WIqxF4V4LYo7n6TqGp9ieXSk48VUPPyBKYfnlW5b
iHnBJA8S/u35EZgAMcgcgy/qxqEiHP/5Sm4f7CG0uOwGO8Vmec76Ot/KFAhZRIZ7
J/lxWWSQlRi6l0jYMGNsNNe3Zu5O1sPOwxKpX9LphaPRY4B1/YYTEmABnP7krl0J
w7gfOAtNZf1pUHXwYE4sn/cAUWz5BdXat9H0aB2YdsUiWpmjAd5O9DvpadZUifdd
ygE9oJrVGz+NKFW4lM8iTBbjGoo3vcmJHTSh9YuCweVje1/Pn795fHyQsLXFFekY
/aqrUdENUSEmkH/Io5tX+irtCuuNoTuEu/KzHTjzHXYrLpK/g3IlhCv1ShsqjaK7
TRRyTMXBmBEujl9A8dKKoLiAjlwN4sznP8uYtckqNRc13k8XRoEkBn+AlxO1LI2d
BzL70wxeVSX8tFTIRgMOoBTEJoHaqUg4Cf7keaieqiD0ds809NQ7AOZgXlbKLjHh
xBhbNG5URjhel+J+TCocb/K1cuZGy5XEImNQazUa3aO0mF1KluGztahgMKFb5ibZ
BEy7YkeP6qiRTNeFf9hxNMS7KszH4Jzin+/B8s0xhWx+MMniRVCehSyM9PX3m4GE
ogUgNw2vVFLCCc14jIRyFPnFORoEfzdztA+/h7UX/ARd23eR7k+3C1t34Vt6OtUu
0VMPdYPPRZNYsPgvZBqhkaLSHqj0lJyHE+Kq1sjHycVvjif3DM4KYzrjMtjE3RuN
dNsE79eRtdemb/aKQd0gIAYh69Lky2pS/3Qajm2Wr84IRr5Y6RoqW1DEPmvP2J41
maYymZRv60f5T+q8nX4uxNc82hgU+FFKJ7gqs9RqEnsppG5b+ILjfZHQR34+JkJF
OLAd75J8BhX6rTj+Vq4zCKUFMd5dp50StLhqB2e9F8tDUe0g9U/9SgeST60imPwr
L2kAZ+1uODweqACJJ9vQ/6FR9l/Aqti9wWRmCT2g1CQLoWrQu/gL9tBNvJiXLKqO
uHE6+rc//x+zF3XoxYIE3hw3Vl2/9QQ4hA1SM6Zf9F9lL6GOeAvimJGwh6x5Oigy
5IdJeMWjAhwyRx/KPgbiLqaSNI2AkzzMAw4ugyvi81+O92R6uZe12KnlBkCND5DM
LkzKrv32YfVqu0JHWbRFAEyW/DDQslakjspS2hp5nyi2PJG8E/7m71/ZAPjBKEor
Al+mMCLtnseac6/nchs8wGmz+QJHbT08rpuG2tSpUowdpsgbOhWAkZ7agaAIZYnc
8//Txoz3965ZD4NJF9EbqxrwczSpm/bf7gpzMLS7enQf1kJA+ikHQOiv4Cb8N9kG
zC1wrRETorySgXYYJ3gP+nzzQtf5Yj5jUFrQrqPObCF1Ru2sTYU3Ky0lRnyNv+d0
GK0TeymZBBUSNjfBkBUzqxQQWFzDN7L1HwIleco+XQgahWHfqu2XOgYtzSVFqAGB
GbS+3+vNLs4IJpCq0e8MTN0saTlx8T0bUuZPNw5wMVaIw75Z+yA/Ih1IAa0nhTiy
pv6jRpQyHFghDM2QhnNl8+e5NxhRBQjWvgHYr3p5vzwHK7iBgyV+1UCZQTbrmb0p
C1dDP15fCnAqXb6osl2TIM4uZOVONI83qB4I0VV3/UYFmdGBN1v94xvu2H5MvULJ
l/D2a3t4yUTfqwNfomb1TieVTt43y8ahLrRsg3BYXsCN23uVRRy1JL2ATr4jIcmd
Ot+AcdgfaCzStVSYijZJ2+KF+pHnxmagF6sdFAa5lglv07ZrZ2a2IBynqGxSuCXh
HHbrEj4hUbysg3KUAnJOyab2Xt9RzxR5EtzHg9L8jT8xWlRadlXfcjRRq9kb7T6B
tnz4NZOOUmWLIKE9ENliCeNTMhqilgjjz+5uFlVd33kGhu3PtmgloJEhqATLjaII
8KF9aVWuDIPLlrCJgqH/UTSYIQ5VAzoslxdp7lcSU3Pkr8et6lXWzeNqKlUuNycD
YW4IBsxBRJue2U5EUmiah8NAHxJxunPgEBBeagbvLj0mxbdaZAKMJWnHr2dLfrPZ
Ez4S3d/3PFKF4Fs/6+Cq03YjBL9onE6xr0LfVKoaFeO3Xw6ym7kTK0tJo4veHRmz
1mCjHPTh8FEeC15BZP+lrZW9fDEFfCyq+/AJSJBJ+yT/LxeVqVaR024AoXRMBGkM
rlfNDxTrOf5GHkoYpv5eficKoPAskC0orbGD8txRT5bYNCHd23CcaA8alpEe5AYv
aYUibqyx720hg9PifWQ1KaTzf1lIVoQox6pGyQIiuF53+FXwwmj6K4oqXqEiccS0
SGbyTG3h0TGcK3qnbkWnH9nCcWoSQ2H2uIKbzWDzKScJm++C/kPPbuSp4hsE9bTv
uxo4VEbwwnhbmu2z+WOxTwIdwiALsAnEzSbmvfAT/ft/Fx5Er01EcvrJpijkNhWq
rCflGE56a+7DahoHVPdCZLif0bO3Zmz6RVQDk7lnwSX89i9gFGg4nbAaHwsCOj42
60gG3gXMzGS5lDLxoTNjWe5Klrgs9rdj1MrgzU5BFyPkVKGQ7dXTj0t/FQDoOQ6p
MTPebvAdlnpr+KACipnbEtSwu7hqT6CCbaEScYkKcCGFFS032CexxRc+yFu5h+9d
GIPSHFVLQphBXiGZQYYIlp0C3ok+0KPFP7WKh+qcDxicdRD4y+nwAkfzvr78UKYp
TtPanAMRUI73MUNuh3JFZEQXP7mz2PaQfsIVaiZbPGIwisZ+Q5AcD46XZG/LuPyA
rpnunyZ2EBu4eTkEbjtUyZrvFi2j14YO41JXTF/Ul2ZQ7x2aGpc4Tk2ohm68sKK2
HJG7dpaHrKAPpReuRPFly1baGGTiW7kdqaIUhOCCmvU+TfFoaJcmkg1zlZ156c9k
H98P+h2Y1F3O4/vDSiUe+RumQQFpM9l718a7PHvPjDmD/WyyA13pIxYQtyoXxA0J
I14kQWzvNNABIuvvqYsh+8378Uu8nmD/ZUHj3xycNPqkTZ8LGizKJWyaSoCOWtpO
AQqnWnTmW7htnTnTJCC/yXAqTvghQ7NWWf0nysuK6r6vwkS4NFVlARja24OaIoqI
543qdzn95vvIq59KAzLlk2p75Wfj4d8IObU28PkvLItgHBlrtZRkb01RZohDOn8g
pCvJNiPSfT5akMp7sgCAMsZOYyWgE8amNSRjlhUqoRxq5W0X2Ya784xtkuMyINIq
+q1Jnr5NesMWmtuyRXq6iMJ0z7+9bItWks+0N0qi/GW8wuZ+nkexV/ldB5lk6GgR
9XVySLmbDEk6ISzHln/KIQ7J0U5IvoWfW3ECt45xrRG/CTc1jzZe7w9K212zpGMU
t/wEuVCsgB0fsXmt0jskeUZj5s9rogYIMCAetckO2gDNnLIaT7SKrIwkqrtnYUZA
94YFksRsg5X1TqAFEKsNy79kvfR4c0vdmewXD1BcvI+85GGzl4Vc4nC1NzFK68ks
qzlI+WeXIsifZLxG2Crki6oyQC9l+lAS9tDEF12GNnkWUz9/lb52cU759bIOOiB+
kAp/PTPD+dl/cQ2+sWlvPLPm4AtM/qTEljDnGw48TDWyKIyGeQrwL/AwfTbeP4hq
neqT3ixsemdpo6+Wfr521Stz5KgyLVFWbD1GFGGXRY03uNegHBMvB0xMxHr0DF6F
BHHzLYBICPipLdxUO+QT9piVi34bT9hUNydVheIjPyNW51BmSEM6fOqv9r2T5f4q
mZy6v/Ngm33Da+He54hnbctgssqDSnbm2WCyWJTS+qYgAH4pL5r4SOXoi5I3s76t
zZp5lS1Ww9rqKrQrj8g3sxury2k1spcUzMO8oXtB9IpWxzUofIkKsArjW+3AnbeX
ye8rLVEFk/RmfcC69dLL/O8yOm5A+LCCuXjJM8+/I3pLslPjBnTWzgYK+29HRyaR
K1DwoAEv/Ky8IpTQp+hCFy3lCduwwfgyqjm6RkxNNIaMGGTy6O1Be6U1ZIAO6pa8
Sc8NV+3iuYRFqA7PZDnQE3N2uJMYKhsdbkV0bUyA6EBXrKjEDL6LICI44qnWZvFi
YQC477/DWHXsgOjFap8CBMqsrF8fMHweK/6Mggb4YC3ZGhKs0dXchcGNgCZTsoEG
idxJK9Fb9po+dYaigD907C33yZpMfqHahIBfpN0xlDwh00ie1NlYLDe3AawrQaad
6RWn1Fizn9H66yf/MIwcqU7PytOfqV/KkgaWSIzj9U1yey37iMem9HBwzXkzt0h1
nis8hoBY8AsoQiWtO2KTz8xbo3T97xY0/JkPytXeNjh0VEp9wtlRCZZkZBo7sBPm
pv/04kB+JeoslylMynFEA5a0a775mZ4ijqkOWgHPvlssERS51Rm0rnx9SB8E96MR
67PTVKnAQLpKuXXHKUYAYUjp5qKSXG7zQE0iDiHnnMD2upVM9U7tDbz/XhkDnfOz
J5Dnn8co8/oqfRnJpw7rh8eoOUwCB875iJcT+enkync5ftbeGSYLRUb6gyh8ONqM
aKnLBOuFwCsehQ238w7qTbg4SanYlj3Oc20PkYdEaxrk9wGveaGGvoyZJory+h0X
CATFesWPhuqbL1I+ZQg1ofI3Tl6s0GsbXwcVNkD/oXE/1uhCEpK/2IMhMM7DhFEO
cwVOHhzjmlVnoKzrbyj2cWyCFXuNQ62TK8Atz8WkH1/CwPJWP+GmouH2v1A4jshX
0MF8yPm+KESuxPemkj9BBoRfRJnfyP3+bKspPWuIdtqXwgjD7pRpWNry8Q+1gbyn
A2tGdSffF6WUY/5rYF1KFLopBUgoGpDXRQF1wI+rMvkYFmqID54OyTjskjxVUCrl
jNkBKSlRpFKN+/dTZUJXia1ywVYjjjnSrPF18PLMfAulOvkmhyBzH1LOL9hiKDjn
qR3eTM3fmA/JJi8FtzPVPtYJyETW6uDfX6r5qAKbuxMDxIul0WPE0MZrAf0cUWuB
9oNqggQ/NlotY5CLLneg321NhpBsynGeNWc/5fyptPugKwomag5iC/dVn0hSWK9o
tlxnrOHt/kQdDg4COlWvHzLDSqcmTgEkEjJI03y54CzwdDOp3CbWYc3UZHFmEPZC
dRJP3N4z1yNGGbDjdXaeNJ9fDGEV8qb6zFzD9dk9ynwcxSPJsD705NtgHWVSUTAQ
GE9NVIRlCS1qUDZTMce2Gy/+nCnKdCMhOqeXXE69bpymbIQM73HLihR0WELRLhDx
+T5k9C26SDB4TcwCAAgWMVoc19eUPQ42hH8QhAaFTc/cFkx7+/JekuzplMESKw3Z
pGnuseMQN3ArkOddMVea4U4jw095qxWHv67i3WT9e4njwq7Bh2SPDsdWvptK66QS
S6RlmOheU82HCyqVLA0L1T5nNwN2QHwOwxE/nZ8FJUgbeDWBLg4D9E81Oc6RbZsu
VHfDmYWm0EUQxdpUMiudX1k0u7AjBFsaodzRMaf6Z2K4g+qbKluMIk5BUpsbXu0e
nwMDI6p35KzWZJKXyxW0ZNJjrmIURSfS9dTQXhMjSMWHoS88tBW5o+p2srAtfrvE
Y1zlbakugyd86hZlAESEvqJf54EXY1+MGr7LOfx3gSrn4NypCZOumWBXgYNloBsO
42dh3//wH56WSJWX3uYpMFyrk1lmdSSqdthtvD2nmavjku1RmcWgAf3BHJTSRPM6
igkJTi3CRE6ZWFjJuyYeBTIPjO3WDWyvvksRr5PqAh8ceO0grAo8NzHwWMRpLsZz
ozeDLCJaw1MEkpPKvwkZ9N4/xgqORvYdxMEZpXIg0o61aQ7qPiLe8UjuPcgDYvs3
iDgicTYgyAHUB8fp8Nwo/ty5iPDtX9olP+b4BeVuPz68qKgW8jcu/pa5JHVfx2U+
GrPFEkFFUcPjUoIQzrfXL6Nl7I7IgxfwLPEZ8QFinyPtRaXSfxHVGPzSOzof7Hj9
WNO18qzgzdpt1O5y+klT2QXqElCqocAgwUueozCRcERtZ1ahkHt43CkMtMInGJzF
kOve8A0zPWioDfZN6Un/d9GjN7oDfqCLPj1Ljxj1jtAeL5SDbDN4geKWD6KYndqQ
lD1TNR3/lSOVT4/Idm8BW3++ssaDiKkJOJTLF/izi6Y+au8socwZtSqkgxRT1ngK
ZmuUWQF+JNdfj7u+/bAK3NBJTryXq4Q/HDB1n8WFrcw8uJ1VUqjXhOtq15NUAgu1
J7FHt0lWt2hoWiPxKjc+0l+NzfdvMd4+tjo0d9LDTL1KZjr034wBpY7/u1XU/XzI
jeDP2jJwbq6OYc9+uOERNv5UZXgWeDQGytk68Ea+gHYEhpzzjDPScF62TeCZzzcE
F83ox6qAZgpTwl/T6bHrXDIDHDNuk+/SqO7vFMkxkCBry4K18SRH+1UTLZH2k4qz
bUooFteDZy7caARV86WjQp+tmHPwttVFUK8cYBdiO/HLjvrznEhnsIq7xA9ulIZH
Ot88hyx0aVigY8fvf4CqcIca1w2EL/EffcgS6Wmk3FwWTNstlygG3ELt2zKm1qzK
ZgZnkKVLueSY21Ji+10vJg7eM0GoOfK0olHwYf/C7O2b31k27AnTFPSBgLzzI9q1
yIk7HLPniQ5QsEpPsZ9QVZEk08w5AUYApBOxKiNmmwvpzRjigxc2AC67G566Hbj3
uJ6s8zfPfAGPawiXF04xaN1ZOF3EZL4VKfjZ6+FP+jCMD1xnR6yzZZ7DEBmdnqDd
71vter5C16wFqdNq+mZZhBELLrt/LET26HK4W2cEjg8A/pmAN8g5q/Ioub4kj+R4
k1jKQHiCJczXN/bKAOPUag+/sfKg8YP2FTJI0M9VGxmoLCxiW9zKS4HIIlvKJ5FC
nl66PIG44aW2P+7bLG+tGq77sRkigfez05Z1KyIcDJht8o5eFarr6Rpzm6enJHm2
Ye9npyFaFybjItFEgu9JiUjfLEWkVQC3FRljYY72nlmYdRHJIkzYlV33ZbYHfJPA
NoBWB5JOvNxbYBymTtGU4vdgag1i73AfoAGr2RYHC5ICXBjVGcO6fZxgrrcWTvyg
Avgue7eaDGJvEnOfhu4iDK7mvvb6dcv8GKFzttsFF8jHekzHbjkMJJmeWOqrHCDh
vJuhy98t9QGr/6rU1i+Js03wv1P4Z4yK/+YTN6o+ny32ah2sHxltTbTQo1BBxXv2
7N2e5g6BCohLJJQr14TSIfxWP5Pok4RK7ZtCbHXsys+g9rcVVi3JN49q4xfVXNoD
KVX6qmctPZbDUQ48OAnn6Faol+ZdwdYcUY0pnIvYoQGvjTg5wg0qfASsIA+rXrhG
6PeAzaq1YM6XzPcZhPniPaJNF3Inpq6PXBP7ancbbFBIYfeUSF5JoHFOY/HWiLma
xxe3sfMj+SZ9BSa+ypsT6X8rnifqWH8N9z0qjMZfxzBKsUAgj7SVy3XmUp7AXwLr
eM/o4XXwxkXTEGJ8NTpwPNKa9CtDfuqvj3POAW7eJfAZN8o4AR0RnKfEQxqb5RRp
gVk8aKCe9drldkosrW83A3BkBucDDY2QZGzUvyPheyJ8G6Ra5osso1UuyRFKLBmu
8wiW6rasucuUTefEnGNQLg9AKfnBIyqn5G7eQxe+go+rmnUPm3dT/+4VH13JYzPV
nOjssCSqDuESVAj+ie6i3hvGjv9feqF5zcO9LRuTf5yAZW6YO5XQd04QM5hAyGum
iy33b8TaY7QQnIS7tk6Phmcs1X9mtLaC8xajgWAmDPZNpSeRABN9w3KPAQKI9v07
9DwwQxGo3KpgGI4SdspXW08BWFyrboHIJliL89Y2A+f7dCCzO2dS1bnPxnD/DYIR
Wb5yyXUAekAGCJID2HzzvZHwpA46wnC4/DaSJPJSzdd7f66tGIdhbWHDKwKkVDLs
tU4AVDiDeIjTZCet8HqcsWhChrgkB9OhzhXAL6egY/x7B8eLPZNlhfWJwy0LVfxt
OBWsU8x4z3uDBGxXs7SM7DIzxGR3bnQPXK+ibUjGU2lmNUbcX8+oLXnEdns0eG9q
UPidjErQWAKpCNwKgpc4YucftOiD1966PWMxxhZXaOinCFcwBP/ZfnzKv7UAdpWd
W75WT1BDzs1fzWdGueGkDM5VvvsBWOpI2MFT9BMM0MYsOAqaP610wjnq+HluOLpR
8dkxqmxFuhTdMww1nK95n3dBRpFZgxKPXV6dE1NXNikiYysjiwHkyRcJw/epF2y6
9JGFIg01WOoFww8e84KXmNWV/hMCg54jF8i+RS1snFSwhQrpOLP3Q3IQFSGl3qBd
G6bMQ+XeF8uaxbNCf0MnJo6LxJG78bn+LwAChcDp8GEHG3OG9n4o8mvYy35XePPS
9xhEdrMJNYUEtSU2+q8gLRbH7kOmhRsfAAjJOoWpQciMIYOwEbpMONNy62PE7NMR
jIaCWPPaHG/jyLOBl8ARXFCjte+/NY7aFW245euSOXlVN9A7wlogtKehfmPsUQEq
IJglkuT20X3TJnwHyyYQ0opWK4r6u0tmZWgDPd9IdoQVgal3GE4QwjjB2NrRPBZi
hkFwKKrQIsOqzpYwhSIij0yekxOxRt5NaHqa450UNCN50Bh6QRAk1hJj1sBbNMEh
KUT0CtEwpRMUNqv2+Xnq3Z9YXgtRj47uoCaOGYP2WAg3wjYounNNcHEbNudsd0qZ
ehU/ugdlRyLdKccdKEZW7B4YpzD1P2qYQFv9jpDERhTL+0GdLoYDLUMNmF3NqwgX
guDIccN0/f9h09jKPCru4Qd1XH9XyVPGjAXJ76P8EogcSU5xoP5Lp3AMzktqHVCC
zxxa+GcJXwcr7X97K/dOYiYRY7T+x9FGiXfcNpzhHf99vpzybMQL/TAYX/M3umzm
vSdFgAqhVoWuY+Nre5V6gz6pEKA+wKdLhA+oLINTIYwE/lskUVEPIlS9GVw3X6qF
/L7yAbUyEqbGlC024gvig/NZgMTUacZNhuvpN6xHTRYU8PZB+LDCjGORXATDwYpo
ldBKUbyYKzBfgfv3ggTYCRnFphqjy5MibnGtOP+/VZIIzDal390+gytM/Ew+Yugb
noHG9RwdLbeVkijxG2FQg7G4rUHsUX+f7Fod6RZBehnafcN7B4O2lKK7fmTFSr6u
sDzBt2xpudLokWZpGlmfDFGSXSgj/JaMqhp8z5L0Y/9PFMQ6gmbNwsPaS6vFutXB
FwpZ2ihlSfCXGU+RoXPgp0yNa57ctcK3qf3B99fHV9bAGLEHF9o7LJ2aFmrjoihN
USdGXfkV2+rNDEZx79TzHFTEQvPtFHrEtJ8bRUYaaAEAUnFDcTKSFwLu858TkDgp
Ow1ExFuGgVK1BzqvMGrGRyUKJ7QXVBmbZfb4RCmFa3k5ltxSzpcT8UDler0gbxop
IzrQLFaY8LG2T1gif6GLl23SY+7JhH8+LmZ7uM+UU59gukRKHp6CkF0bkY6rbM30
buhc5WVkuZtjTzi85W64fHp6Aj+Y86udwmVdHJ6xdUzK0d7HVMy00bC9gpZtl5k8
zhf8oTVlAv+JhfJvGR1EBaPV1DTLheK5/+pd5s5Vprq1omcAnRhpulww/mZrSUn8
gWzSxoqQIsb9LWs23xAkNK/hoNR1L/9I8/vPFcqFDlcqwLOxYN/5Ks8rf0wzavPk
hmSGs5o46LuaUmqNDs0P7TaMi+HKLIVn7fQ33IulVS81BR8AJ/GMYE5X+vyss7c1
vy6g15ZVfTlZewq3GwLpZUHkuYDygFM3vGQMPUdh/rWM04UZg6rFhH9JVT4RVOut
mh537ZyjB6a5xv7BDquHVGqbJ5XLAfuqukQeck5dDHOpijV+gOZanByFIibLhj1r
q2SL7PGEvVgsBoE4Ib1z3TRorM1/ePR7+2ovqk2SbYXCIRq9IHzSxXdRh1CsTJrj
QsbeABBjKAR7mINytJNFiFWB+VvCCFe6C8qxscPeFTOw5nQIbwrO448rMFNX6e3h
lV0pIkX0V5pfTSZ+Y6HFgWDbYQfXFEZISKWuMx4NVznvdXs+37ZsecHTqsH1xvl5
2Hp10c2fy7XdQZgIktoJqleF5ovOjdScsUyoAgNGe/0ZOW0DILEDXx4bRqwllSI5
U9BibCmcyEZ6n1Ha27oJbGq4O5jpPrdodqUI2jC+u8YQ/h9ehdcjm/1UO4JhmVzt
oQ+nMQQ+HOlaESMp1AUZHfRUTxd9ljdu5hrAezb00+KNLt/9VcISd7yXUBt9iSv4
HJ/V1rMQ+fB1+XIBtL1NoUrHBvCHbVEIx/8xGpZMtzwDSt9Jua7IrxU1ioEcu0S0
7JsmJx2NfWexNcFYOE+aRDKz0ACFOVjYy64GLOseebQP826dvlEBTIzd3VGYikn5
XYcpHYY59OtjWz+E5UEJi8aXbdxq33IbF2tveKCkncoOxdV88pmdX9zivxZtX05h
RW2Q2iHKwFxrLRff3wI6d9kiHbXKsABs+LOwVziOx/a/xq7P8RQYUlO0jA7dEBcN
M0YzYgHDDzWOK3RpjRTtxc0hdMCUWQkJz2C3tLberUpeSYBktRnjjRQdVFFycxzB
ctZ/isM6B8GR+F2XaLgP59aQmya7lqaYxU3Oefvf/RbAbLVmbHOzJgd+qr1iHtP2
PMXzwtypsKunsDb9XS9xv6NtLAVBBXFp5EEbWEFAFbiq1S84XuUkM3TVBfkxFYEM
/5dcJ78JhB7a2KF0zcUomOcLuUnNiCWxvCwwuabTVd50MtxB5GhSAOVhwfBZOY60
+mEEF/rFZEhAy5XY8cXh/w8DAQDBlK4B0zqjJF58x5WwknHEk07GZoD/Dv+A9ayA
XOMYrIIe6o/LAmKEFmS9oGg0wZyQgNjPxJnGPoRVlUutmxgHE6fGTnBHL6v6fByN
3/lkEFpqPlKYuwMwjynZDxsP0dMKv+9mVsXERRUvdOjCoopO8rqYXnOu14oFD3kr
8xsOLHneczGOZvAllbvwuSL+2XUh8ZkVX65A70+AR7juiUx/nQ0VqI+MfSD3S7YC
07v4T1f1r3kPUumAlNvJd8Za/bbxLB03Edizc4A2c4w9AtnS2Na+TUuZ/YKeEqAk
1nQbqAWZOXDvv1aUlSC9jFThEqsoxrJTnVtZD/G4OtK+kjMs9knSCoMWTGyH9SKB
5dwKzQ8t3dzUliQ6//Qi936eFRn0dfFPrDVmduAK4Aj1igbg2azoBYPtTHqpZ99t
9Py6NZRyXJAel0Mf9LGxSZzC6SMvg9hVx0gl2FMdCOtf+drBEFsTJIvO+VUbEcMZ
gW3p0U/9T27+P3AwuzMnGZGD8PaHj8wGSAIn20Y4C0eCcLgowAP08uY0jz8HN+kP
BhP7F9f9vwaFoKYCYkin6Uqrye8Vpl4KdTKgN4fvIcWpbb59IhT7JJXLJAziRNhr
zEzPGkz8cizbqMCZA4xfm2u4bNeQ6tfDKtDT6GJSOrucPGKRfYM/Fm1BDsZpTmON
rwmGeYQW53AtMEIBKziadwg/6G35j/oVsrxW9sh+76wr079QkMmwDUX0kCeROUjn
SNkqng7MfAoqbv+x+yDqQwHFXQNg5/xJ2Anb8yCqbq1sXc67R2z+bqpu9esD7nxm
70OowCopawAMf4wQMFAb8eI5q6tNgM1sD48jZVOu9bp3qIO8opL3cHtoWS2qnWpg
ZHLYWAGBNN/WgOhOIiVHCmc8/8H9JLaa4ogWlJmxoxv+nXHQRtRVOqbI5VmqUZol
PMiw1L0gAR/JKmYU5bclQC6mT8L+vBqbdVuxC/td8afjuGhJVlGShdeKYB62SMI3
ZocYz47rFEqMG0d0BI93G0ypV4Bt5tOeXChLsddDgVsJ6KpEYYzkesVxrqWS+9hv
MLHcSJtjADw95+EmjsuqMvF//qMLA/NvXNN8Utlqea1yhckTQkCJ3DB7dMirK8YE
8HFAbSCGEZ8LnQ51pVbiuDmN0sS8Jh9R2T4C08CxACOZ4kmgyWEnGWnK8+f14AZg
Z43SOXtIdJWwnTZaz/SuCNfSJzVbu0sXjSf4N/5LrkSeI/cQ5YBC0AFMS1ForJHz
qQNW/L4e0IEiJuSodVFV88b7A1wJOKeMX+WtytTLuegPz4EP3og+9yVVM29k6beD
CdrrEQacWitiq+qyCKpyNdmvyaLLXucQhLjSMrrx0xkU1EagEz/puG+kggV1OMWJ
rV76BiPiirH8njjBX4bZvJH/PzxzUBdkHnO442V6POdtUGtw9OVqzhyfMnurM0Ug
8WG1WwysxPAXcz1YESEyfrNjpQJ5DN7MNQSpkS28a1yGrXQmyBaTWlwbga+8r7id
gVOb9QEe11n4pdkkJG8m4/T5zZLgj1hgHACisjNZf0kmsCBLx1btwBoUkbxKbQG8
v5GH+KdDGmW9i29ZRySYL/0zbAyhWXd662X5xCO2P95h4SW5KD8gqp68mx39VffI
AxwEb/ex96JkeYIQoZ+BwE+OXYM12UAw/m9IeiXGIVl9mnoEUkmpjzfuQN0gS7+u
vl6KAq8HZ0gx7GCYIC7fvItKlURTc9yuMn+nG5XOfwh0G5vJddloSZ2KkEyzR5Si
oq8Qi2op+pBUBmZXKBpNq5m7zOxdXbtv5UyFc1JHhS4a6L8ysoXcfeYSj6Cbx3js
C6IT3IoZE70fkZGmQiu45zNGSpUbTMRmupZwH9GNnqJtBjcRQEemUrWooie0Q5vT
f6jASYva4TGIRywIM9f3jz8+fgAAP4RS+OKihbyUJnm5pIa2yMT825QCEVnC4kXD
frA//6OXCCAsLatp9vTbG+WL+Itm3JejJyZbd5BIXfmrSyiUK7fjvuig6l83cfbQ
saQpNnnXG10fNmqRPf4NvAUPn/22CxaPcCQN6CpZqWxiNKvgUhLlBdnsiCZv86eI
IRNtuJ4ep+FUVqZ7oCE2HWAc138y+ZoCyC+4aCT15sD8n+9sz776UfF69QV6YhqD
C21RLcnOLG+T9NVbyLCe9ueiI3jy4qhRPw2+BCc47kWDHzEw1uPX/bJSxwwS1S0r
x8vTyoOTqSiaNJudOPd1CDJ+DYHEQaOeZ9Bq13d65WSCvIAaw8JWiMZN4mZKNSbf
ubst7eavzEpmLUCR9a6ahsVlgkxa6PPiZvrE2GXe4qjTpzFRgYzus1AOyHEiiB4c
l1NZENNRrIGz3ZqRTfnSwAEjqP5DAJhXVYibgbkt1rnj1tW2m1IY/WF59JVvwDYj
xNqIMnlipO0MzxCjpHNdIYwylLyyPYXJMxJAheVDR3QDbhnk14XfkKPqwJnexGkP
kyfxfuI5fMuWAYAicdWCGzle7di4i0JvMtI/TIR+FR7dDHoMg6dHuyBLxXbzJ1LV
TA/6LIOXUhjnRU+3TvYbwk9EN3oV+bLQMB6BJ+l0kCABKCBKqX4NR1vw8tfQhcyP
pMeuVMuiTwdogcao6j5BhJ4NFqIrHTpgisfeCeDmvqf6Zi8/0T9dha7HrGrlqdJR
0G3lKAKjRsUfzNkASCWXI/We02q0d9G68KO0mKjR5RE+5qGE4NEKTFsrdMMIfwxD
dBFp38JHk/+pTga88AigkHgxb9y4JwFSQzRCwk740S+X7xFbC8wa1/e6YsTbmqsN
Fr4gxCAaeZGqiWxnZNbwfPweM04uQ4vv4SV2nbn1jkI7IaPMSPm7BiGaLBdFvShH
dSK9TyRm4Bh43ca9uyeAcI+OPzUdZTRRWWrvqYZLKMLDQna30JGdNbpDCvRxPFmj
XCbZxhXUGabz1C131oRBpUPN0OFwMfeCTKnQ+vlPA8/45s/kbJ1Y+IEy+F2lCRi1
Xvlfb7qEXtwaQAfPBOKiMxKYVfi299i+PjMks7BKtZFLT3Jru/LkdE51AFPAvhnG
xl5qCzEUx7EjRPAG7Kb+aP1RExquROKV1+2EVIaJdnb8F5hS7NmIYgozAaWUTSST
RdXKSKmqA/ZNxI7Rmu658U2PTGhr+OxTu3jRwICn0/d38hgPHFGIJgjHueb3tWZC
ERyOYmpw+3Rucd97RCbe2oTAnNWZ92S4sZuiQ5He643ABIqkjtAKpB5+G9dPS9Dz
U1EimNIR02bwmgsuky8RA4M9/cuGRxllANz9RjfmHPkn32PtLK5ldTG+Frpkrvd9
4WP3rnPua8uC1gmSt/9fvR4ujWO3q6x9CP8+UWFiOGGcAncdRBdp47rxHfPngXaL
ATjA2wj0o2i3uGBYpwREO9Rj4K0Nei3f65GvXW6YzQkt4MgiPBH2pyjjmt463gao
ATrTGPuSu5yAR/2FzabLFe/LPAX48PZ27jWJGfe9RJSCFliWPmICn5bqZk9azWez
5ESO7uXGbjaMLhMCjF0GHXoyxNeaFD876E858kpuP46JA8UDhV9R/t72AhOPq4Hj
gBiixhS4Q+6yW6V/4FP/ZMB9KhPmZLMrBN3jMinwJaBNVI9soODzTEVmHB6HFUrU
6Q9MwnTVFOUzaB7uegXuEdgZIgRajw+wTe0uXDx6/B+ZF9a6/R12+2/43HjWJzbf
vhvdyg0eF3mOwSFPpSsIi8vD/97SKvC/U8cypw196Jkb0L+zqEslgInU5T8kNpM9
N7HO1bb9FN3sc9Os9dfwzzOeO5pTMlkLy6S7tEEqfwkoZPLWEdgwuWrgCeH8dnQn
Pw4EVePlf01fNYJUDDJ8gVTsa5jdfIsuzo9xTJ9xhhb+JEBmYebiO1ZjvspVpKec
pyIHM3cj/hmpLm1mg4BOn409XuNrZm5S+9ExFQ01SfyQQHDJygkQ2OgKwvexQ3Si
49mBVt4oyPRer9VGPjYjx8fXUa8EILrce1L9j+bCCBTtNkFtb55zux/P228DptHl
BXPACmcv442r0KhoDA2nU170wiXPK27p4nh7jdn4Xljh0TGNBBjxEjPt6bTJm6Ih
EFYE/IzjhoalZbOlS4Yqe1GHDwjKioHEPhivqZc8Ex+Q+eZhpiJDZw/FbgB2KU9g
O7hhiVBBXhYX0mAM7uobKufZIFX1ukvbpypkvcSO0mC7IjcwU/GXpRil5dhzAQxu
LOCi0DwzIVnyzOxGPdaAEL8E92SnayyqjtbZ/sieLewD7ZpS4op1A7ccTuxrhGhY
Cl33YSZ0EHqYNimKyDRYC326r+FePEeSc+m0YQE1pxcTVY9C5hybnv/QfMqUm3h7
k5kMTOOwj7Xw7oBfb1T9Mj5fhtqsuYcg+eb2qaX8cirv2UoXGpYiYP+H6NcCcGwG
drPrQH1cBBgzzF+4LTgHwgxF902JjClgn3NjcB5iX9xmNvQ4U3xARXRyB3oI6jf1
nQ0T9lZe/y3GHI1tge1PcwDJpq1+jJhBojgX2G6r4OTuLyeszvGXBeDdqc4KDCCj
0CLUpxd3rQ6H9d3YXe0LhZ3fjhQS4xxca7rbvcDFx91yLa+zxF/YQtYFSJ54eKzS
m4yKAFyqn0ensoHHFerVjnPbaqeVzPUYtc/qGjFC2iUfvKl3mO6dSF3TDm7rA0XJ
J5oroIN0RSG6hxjDg5i8z6pLzxAsAbTHbaVQU4+yDC2QZc+FiK25lJzELzjRSMHM
oaqEgG/PmGBXsuS5nnlYnNi2AAf+xOPl6LmidcpHEH+9ZFKyHligRljpvXPqQgHY
/TZ+at/E9XqrL+u23QJHP5wJh0hns9pPOIasuT2cVnCixF4SPgp2WD9s1GxHTY48
uz1/qUaQ+0vWiGZxJq/Lr0ULMi8cDPD9r5Oam73usIUz4vvwkZBz1AQoJCduG8n3
r5csFsMsDlfLxq5Q5cGzHBX7xWxO1nOIJMEi3RpihWlF+HZ9Oo5Ru9ymSPwoRSYy
ly7KfEVdg7vKQ31Lg6jfJYnCTCfl4WbhUqSaiOu7U7ntNJpB6GryUJCyH8AZUq9c
YhygiiUoH6a3ftKirVHA1DwfKZWxh22QIfeavlq98pA31VNOKFGZ1yhSNmY4U3WT
5+sw7s6tlmlhITggaTDjXyWONGhGcaVOAdSkOmwmBiSnVmCmFIGikeClTiLW5p6N
j7C0oFavgv3el7FIvBmPIhQOf0C07+jJJdufjYD1oAdINHQVU5XQUvjZcjA1Ghfw
qIwlTKr43Z0yWqWmWUPrvyWL5YlYfo0XE2L9zYAUvm0wsP7WJF5Kg9XAYeRxB7sp
ZV3Ze8N0fdYQVQKk78hJFzgttiS4SfBVgtk6lcEs24sxJNgGXrLe+FeQvp6mrxQn
XTASzODlat/oMy2Lec2UzmzD6qKaw45bZdUTvm9cpFtZYT5PjQ8DbdmD2upTcik3
TxI2/3eycZSSQe144Ffd5fHIbGWKYpVH/xkWlo0IwYZZq2WYrLjM5KcpLLZWE7qO
uaSkhKemnU/WiNoyySeS4lO2ZfgEmfjzUKv4p3mL98vkElWhdzM14yNpntqHA/4r
R2N6ODZ47keWzmW8irj+xgnVkr44HZUb5zMeUwAMWz5qTQmHxiR8P2fH6aJO/ehj
Kyv6UmnA1iIAAbxdieruxQk15Ybf6NbeMaUUCMXRXS5U0T00IVJCnHSDxZTcIz68
oGnYK31AE3kvAGTCyLSYkwiBKuHM71UED9HL8HNgtOO0DymDu1MEeD/41qRpAHuk
p54jdCyQLpuhE2JVAEqEWlKKDqFR6Tt2Sk3aI67G9tMD60t6ApSE91RgcRAoD+Na
wCEwJPIW07gzERT2PP2vQ0LhNN8umVr4kGzrqh33c3VWc3VTan7s3p5hma5fajSg
1eg7GOlCn8vY2FzSQu/RO2Vx/53TtbHBHZtYkqhjVq2Dm9CpX5oHXfbPWhLwhP8F
tULG0/W8ac5ezdj8SAjKlx/0lfg+2gCSs9aFcarc7dqlAQilaiujuwNXW1KQ/otV
njfK03v0MikJ9bwvB5zyX2SYJH74HC5LBzKspVjwUsZaMTVNtZl6AvTixL93LGGK
`pragma protect end_protected
