`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nTY63gTfZKtDvGXutDsg4iv5A0vVkNNtJgSdwJkm6IyHM1uvrjWQZPRyx+5d7Rur
v5UWEVqgEobk0ZQETApGwJE6pk0H30PhjegNulB7YdM6xi2x18Io9Ye/1nTqgJuO
9aJnrBPzXrW3gIMge/9L8kyFE7AErTSQyY2ngW5PJuI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3152)
nBEUHTi4FqgTwpJXl/Sgv84POl/34vDRpHyNxSoKT/C1gLA109jNKeWZyHcYoBzJ
+YT0VPPyPIlpftFF+Inbk1ajzP21HDlu+vb84RmSsmyz2NqVL1y89n8gv/9QaFiS
TyoNPH1WJks+Sir7Jhem5XpePbsrm6p7ZzdeFM/lfLkBwXss5Ydw4ZTCUxeM5qbD
mHJu8XYqlrnHvlkdqLEirzW3DdmwkoYN/n1a+dlAKGQeEM8G5yt2LrSpwb+Vp/zI
iR5WCig3YAqmJmknE+2do4Ue/mMsL1E3lyjFaLHQC1UE3GyY+izxiPQIPFF2dGFP
14VPoq/Ia+CWoArr05D1xiVRXMvxZv5Lfe7HbJBTzXv/VrPbfOijBtrF7GayOs1V
/LwU5pu5PRU1a+o1i1cZjYkt3RYHgb/vHrVtoDvAzImd77wmtsCKeWWQdjFdiPpw
THS/LKTPa1PbReVmEcM9u0Mu3ECtKFbU7Eu2IzktiBuBPDjc8uqHAHzaXZK6x5dn
k6z4sszlh2dLyjMXtNfBLFTc2RGh77o/k9CmMlKTTs2uOckWjmDr+Wgbbc9+Pi6s
OwY07MVecCJqVYgcdJ93e3RmmpgHuee5OGKo86YBOu7nbgKFdB0ZOi0zPWjwyHks
Xijnra/emTiEWaF7Gs63oG+NBtSu9SDL0iKjdgsf3cyWXko4OCrTxMCIJqTdhZ2R
UliYCRNyz6mtNtpCtnNjdtVQLzTDM7FjlsgEUdLNmsuqqORXN+QMz1li8Ebi37Y2
f6aTkAePilEZ8S0C4X1qsl4h0M5lycsEXCjoKMaFZJv/EOxnx+AEwOMlBqnO378W
v2qMX6z09C8ZpEguHD6EB7DclDkuQyZlgkJyeI5Kh2xtS6V4Etict/RRWCQRaKhq
f0S3qBpqy0MLxYyC+dGg1MiXRNDXGy879wAbiVQ6XsQqViaX1F0RY25uossd8+D9
7LNnrWWYOuHMlF2S3j4XiZvSLXUtrsxBc/cfg7oa7349UrfGu/FQKD8PfIArRC8L
HD5unJSGx/IGTjg06+WuUfjiWytVia3nn5irKFtg+wqI/kydI3K3IyrsebGAxNYx
TfCtdzQL7aTOM/iBRDLo6VKkaLs0LJX4pjo1SYtk2ti6WJmBNh7xWdjoyPOMW0lY
kDtjNTKWTD32VPrdTDDLeVyvCZGkW4ZgLnU3hlmUf1VPWVA0GWpb7zm1SWnkEeqU
pY3ksnpMmlGMHWFI+2/o0zWSc20AXIGO2S3grwaGCgm2SeVXO5kRHPbQpMtIwAM4
i8xPkeDlyMicA/O4W0NI1lnlsARWEfgEbgjC4DqdztlgVzvdl4i2oEseAJ2+/oDj
ayI9Hr8bDnKOON6Db7fYFUVSpHdN+RVcrOKgZkc/qGuw4F7DM43qUzu6u8Ql12yJ
Lingy6MF2vbmYX8Va6F0sCI9X9NjR1WXxnVq7Wxyb+Iogx8+Lko8XhY8drkEr046
Zj2hQijq4FXc9Q9UFJbIKxgpUBrOiW6KnVMow5hDR0iP7TTOW0lsreJX5z4be/qU
lpH67evLyatEhCB4+yBu69zTmhU0CW7APZsTlp0/lIxAI8C6FDtx8bKLGeN9+iqu
Gxaqe9CXdyslUQHY2C8tqTn1+tAoRrZYBSENY/m9ycwcJMwyumjnjf7rq9UIWO46
QVz+I1KwN/K9jEXN7rdmiP1O+JaE9/OKHnTsoy2kBcvshy3DkR4RkSyx2OviRDhM
bvojBjzPTpJeqdEOXKeI9+WR59oJGMGpMzzad0xqaKKOA3SD6etHHtgtnt1+oJNT
dfPQOM6YAxzFRg2EylNL4RSWQRqXJIT34ngicJkT9uMGTrZExrWSHmh2gieiY3kh
o8ezs8amPdmo+aVLpc8qs4CRSkhvVqaIe1wLrYgblQSeKyqROfpCyyIZWgbYw2u1
CNQCVY+/Kbxc+2pv7hvLXXybAAHIonQS3f8i0pq1fobDUUmzouCy1TINVp+UrVAZ
wduNPnCMAD3TAQbRTaWmzLkjkwxjPgrSOg6BAmugFQCD/ZWcHUlXt7kjQ8BynmqA
yjRIIwC5NoUtvR7/+CKBQzlOso606Z5PmhA7zDUYrYwb20LV+FmdfbRd8f9NIJFf
z/DI3YQ9DSyp5CbT52pha+NqALe9sy158kXfzImJhQfZC1D6GjQw2IxYE0GYyp7C
7g6IvtHjXETrspBEYg1gjXARCbrQIiDuR3TmRBdvm6QmmYP+GSFVu/hLBfCRRf4Q
Z6huNemumgbhweaAap/pGRQ66ZjOs96scv/OXIYQ3O/03YkCzuaE1DLriIg+Sb3K
GvMthz8Nz3iGxpbvuEWIlLMVuIwqauNTa60Al44V/oB/9+Km4z0YYvibg5/jDhlk
ivgyyR694mN+IshcAAPcRzQ7pbxK7tJU5pnVyMGpwwBOYM/TCmEs9eSl2ZtJu6iv
Ii06haGZYysAIHKb3HXtPgEyyekA+eDYOoR1jSRzszDiJfVMXcup4eiad7uAy+0i
nR7x+AgU6fa/X0z2pIFZ6eAD02Y7KxytFkIORxrqScyFv/y2j+q6XeMm+L2fcr1T
51xeXmvSMvPUUQVUAfBb0aHBBYY7ZxZCqMeK1vLoEJGqyV+SaR2gwtGWwzYiNOdL
VAKMN1vcVIQ1mO9/D4gV4O55U64TX4pfpIDGaD8dOSNUMcmOho+eWgAD2tOcZ104
yDs7LTgQNz1y1Uz+tGNb2xGuon175liHRC+A/7ipAKls0xjO3UKIuS4oLKYp7dWX
+nKNt3PgrlHOTJO0JNTQKP589qInbNybkt6937KJVOA7cN8XhC4LBfkaC5s4Bor7
eYdTRt9HlzprQPaIKoJvn3gjBd9cfbDC/qYzdWTRSev1/qftsgiGq2PpdJ0nD2BG
Pyyp2Vkdjby3EjEh9UDZ3rxBe6IdbR4DBiS6bu3gXAHL6VGs6B6DWy+uDCe+CgYf
ChNi+4b+p15qOFqoD24tWo0jRjpAllCCY8hkFxPEk3m28mFzU7hk6t1Z11Gv069M
aM7p02gaKXNFgSjx5oY8ntqOdOi4vIQiCyleESx5hSoA2DaMmaWwPUh/zF+Z9TtN
HIRc+QlraEdHTrWlkwLjVtujDt3Slz4VqIhfqcgn0SzG3kJlT5M7Ay7OXnmGqPDL
R/KlvsJRiwXrf/UBeLJTaf13Y53UQUGh8MPpEfhLdymdG28AYS7EfBBH0Y69WdAR
ltRbw7RPcfYeiN+EdzECs6XaYK1es0xQjdPIhJSckUiAKt4mOUJKDZSFFfmGKSuP
ETTN4/uz6jhzxU+0OGZLA7HwTY1U9T0HIVlVD/trQk3DigaXLywNbjmAvCpfBmQ7
BrTWRUesbQ2AHa651iV+fv6v6EZ9FcpDAS2+7teT6qEIzFC4D17ws9PY3s2PS/LX
+QLeYhAsgxj4rvHsa0VAI7B+Z8In3qJVohPt4JPPTHAXjLNqyRHJEee31pEcHof7
soliAckShFtpg5mstgY8GGTTkZ9FO0CvJ03gy49zk4St9ULy16iQYBC7Z3gJJRzI
HEL7bINBZ3EryYAltoC2DBvBs1cHUNCTqWlhy9mXdgjePclxJrwpZdn++JhCB1/q
GAKV2MW8lzG/LdAqT8aIrAm0xd2FASa7NydlR9Trbp9KjWaxkYSocNwfFL6/3xkk
vouKYm1eD4ysI8unvrNkZCz+tPzpMSXC0msqvUl7GG3hntaPX2nFYFnmagLr40Q3
SBVpg9e1zXvLtuUPRuXIYoYbx/qr9F0O9HoTxdlfcoWT4Udusk9Ck8TR4Wzw+vs6
UtJMSVZT6f8s8wS1cRijmmQxyHhiBNiEPOa2K6sU9k74RVpYmUxJjA7DwNs/rOxq
bpcv83lRE8BiviKjkVTz0b553Yg+q6T67csAOGzWZDDKCtSnoLFzrRUwVvG1FR+g
z1NXLnBuazuU8lOjfzPmTE0VDbMZ3VdBj8esiz3UPjBBdAZMBpPmoz0HqUu8T+Bm
ceJZbbi4+VbhIGDyhhWGXjjt1tC2ROHaTltoX+rcGz9GYUPVc2us1J24F0Sta4ny
vTtyp2aOTv4afm1MhlSHAY/+gEZCob6XJ7f4HWAkF6ckyWDEXfdAuGK5g419veu2
evn7Rq0ZoLaBWZjvPCdihnJYAkPBCY14+H7JrVGg0e3APMm+N0cIUU0fChWol1YI
PBsdpv+ykt86LDwUX0zf1tzPhZ4Ib1lE4pJXYJvMbn4=
`pragma protect end_protected
