-- avlm_avls_1x1_tb.vhd

-- Generated using ACDS version 21.1 842

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity avlm_avls_1x1_tb is
end entity avlm_avls_1x1_tb;

architecture rtl of avlm_avls_1x1_tb is
	component avlm_avls_1x1 is
		port (
			clk_clk                                : in  std_logic                     := 'X';             -- clk
			new_component_0_data_in_conduit        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- conduit
			new_component_0_dbg_data_in_conduit    : out std_logic_vector(7 downto 0);                     -- conduit
			new_component_0_dbg_input_en_conduit   : out std_logic;                                        -- conduit
			new_component_0_dbg_output_en_conduit  : out std_logic;                                        -- conduit
			new_component_0_dbg_write_data_conduit : out std_logic_vector(7 downto 0);                     -- conduit
			new_component_0_dbg_write_to_conduit   : out std_logic_vector(31 downto 0);                    -- conduit
			new_component_0_input_en_conduit       : in  std_logic                     := 'X';             -- conduit
			new_component_0_output_en_conduit      : in  std_logic                     := 'X';             -- conduit
			new_component_0_write_to_conduit       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- conduit
			reset_reset_n                          : in  std_logic                     := 'X'              -- reset_n
		);
	end component avlm_avls_1x1;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_conduit_bfm is
		port (
			sig_conduit : out std_logic_vector(7 downto 0)   -- conduit
		);
	end component altera_conduit_bfm;

	component altera_conduit_bfm_0002 is
		port (
			clk         : in std_logic                    := 'X';             -- clk
			sig_conduit : in std_logic_vector(7 downto 0) := (others => 'X'); -- conduit
			reset       : in std_logic                    := 'X'              -- reset
		);
	end component altera_conduit_bfm_0002;

	component altera_conduit_bfm_0003 is
		port (
			clk         : in std_logic                    := 'X';             -- clk
			sig_conduit : in std_logic_vector(0 downto 0) := (others => 'X'); -- conduit
			reset       : in std_logic                    := 'X'              -- reset
		);
	end component altera_conduit_bfm_0003;

	component altera_conduit_bfm_0004 is
		port (
			clk         : in std_logic                     := 'X';             -- clk
			sig_conduit : in std_logic_vector(31 downto 0) := (others => 'X'); -- conduit
			reset       : in std_logic                     := 'X'              -- reset
		);
	end component altera_conduit_bfm_0004;

	component altera_conduit_bfm_0005 is
		port (
			clk         : in  std_logic                    := 'X'; -- clk
			sig_conduit : out std_logic_vector(0 downto 0);        -- conduit
			reset       : in  std_logic                    := 'X'  -- reset
		);
	end component altera_conduit_bfm_0005;

	component altera_conduit_bfm_0006 is
		port (
			clk         : in  std_logic                     := 'X'; -- clk
			sig_conduit : out std_logic_vector(31 downto 0);        -- conduit
			reset       : in  std_logic                     := 'X'  -- reset
		);
	end component altera_conduit_bfm_0006;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal avlm_avls_1x1_inst_clk_bfm_clk_clk                               : std_logic;                     -- avlm_avls_1x1_inst_clk_bfm:clk -> [avlm_avls_1x1_inst:clk_clk, avlm_avls_1x1_inst_new_component_0_dbg_data_in_bfm:clk, avlm_avls_1x1_inst_new_component_0_dbg_input_en_bfm:clk, avlm_avls_1x1_inst_new_component_0_dbg_output_en_bfm:clk, avlm_avls_1x1_inst_new_component_0_dbg_write_data_bfm:clk, avlm_avls_1x1_inst_new_component_0_dbg_write_to_bfm:clk, avlm_avls_1x1_inst_new_component_0_input_en_bfm:clk, avlm_avls_1x1_inst_new_component_0_output_en_bfm:clk, avlm_avls_1x1_inst_new_component_0_write_to_bfm:clk, avlm_avls_1x1_inst_reset_bfm:clk]
	signal avlm_avls_1x1_inst_new_component_0_data_in_bfm_conduit_conduit   : std_logic_vector(7 downto 0);  -- avlm_avls_1x1_inst_new_component_0_data_in_bfm:sig_conduit -> avlm_avls_1x1_inst:new_component_0_data_in_conduit
	signal avlm_avls_1x1_inst_new_component_0_dbg_data_in_conduit           : std_logic_vector(7 downto 0);  -- avlm_avls_1x1_inst:new_component_0_dbg_data_in_conduit -> avlm_avls_1x1_inst_new_component_0_dbg_data_in_bfm:sig_conduit
	signal avlm_avls_1x1_inst_new_component_0_dbg_input_en_conduit          : std_logic;                     -- avlm_avls_1x1_inst:new_component_0_dbg_input_en_conduit -> avlm_avls_1x1_inst_new_component_0_dbg_input_en_bfm:sig_conduit
	signal avlm_avls_1x1_inst_new_component_0_dbg_output_en_conduit         : std_logic;                     -- avlm_avls_1x1_inst:new_component_0_dbg_output_en_conduit -> avlm_avls_1x1_inst_new_component_0_dbg_output_en_bfm:sig_conduit
	signal avlm_avls_1x1_inst_new_component_0_dbg_write_data_conduit        : std_logic_vector(7 downto 0);  -- avlm_avls_1x1_inst:new_component_0_dbg_write_data_conduit -> avlm_avls_1x1_inst_new_component_0_dbg_write_data_bfm:sig_conduit
	signal avlm_avls_1x1_inst_new_component_0_dbg_write_to_conduit          : std_logic_vector(31 downto 0); -- avlm_avls_1x1_inst:new_component_0_dbg_write_to_conduit -> avlm_avls_1x1_inst_new_component_0_dbg_write_to_bfm:sig_conduit
	signal avlm_avls_1x1_inst_new_component_0_input_en_bfm_conduit_conduit  : std_logic_vector(0 downto 0);  -- avlm_avls_1x1_inst_new_component_0_input_en_bfm:sig_conduit -> avlm_avls_1x1_inst:new_component_0_input_en_conduit
	signal avlm_avls_1x1_inst_new_component_0_output_en_bfm_conduit_conduit : std_logic_vector(0 downto 0);  -- avlm_avls_1x1_inst_new_component_0_output_en_bfm:sig_conduit -> avlm_avls_1x1_inst:new_component_0_output_en_conduit
	signal avlm_avls_1x1_inst_new_component_0_write_to_bfm_conduit_conduit  : std_logic_vector(31 downto 0); -- avlm_avls_1x1_inst_new_component_0_write_to_bfm:sig_conduit -> avlm_avls_1x1_inst:new_component_0_write_to_conduit
	signal avlm_avls_1x1_inst_reset_bfm_reset_reset                         : std_logic;                     -- avlm_avls_1x1_inst_reset_bfm:reset -> avlm_avls_1x1_inst:reset_reset_n

begin

	avlm_avls_1x1_inst : component avlm_avls_1x1
		port map (
			clk_clk                                => avlm_avls_1x1_inst_clk_bfm_clk_clk,                                  --                            clk.clk
			new_component_0_data_in_conduit        => avlm_avls_1x1_inst_new_component_0_data_in_bfm_conduit_conduit,      --        new_component_0_data_in.conduit
			new_component_0_dbg_data_in_conduit    => avlm_avls_1x1_inst_new_component_0_dbg_data_in_conduit,              --    new_component_0_dbg_data_in.conduit
			new_component_0_dbg_input_en_conduit   => avlm_avls_1x1_inst_new_component_0_dbg_input_en_conduit,             --   new_component_0_dbg_input_en.conduit
			new_component_0_dbg_output_en_conduit  => avlm_avls_1x1_inst_new_component_0_dbg_output_en_conduit,            --  new_component_0_dbg_output_en.conduit
			new_component_0_dbg_write_data_conduit => avlm_avls_1x1_inst_new_component_0_dbg_write_data_conduit,           -- new_component_0_dbg_write_data.conduit
			new_component_0_dbg_write_to_conduit   => avlm_avls_1x1_inst_new_component_0_dbg_write_to_conduit,             --   new_component_0_dbg_write_to.conduit
			new_component_0_input_en_conduit       => avlm_avls_1x1_inst_new_component_0_input_en_bfm_conduit_conduit(0),  --       new_component_0_input_en.conduit
			new_component_0_output_en_conduit      => avlm_avls_1x1_inst_new_component_0_output_en_bfm_conduit_conduit(0), --      new_component_0_output_en.conduit
			new_component_0_write_to_conduit       => avlm_avls_1x1_inst_new_component_0_write_to_bfm_conduit_conduit,     --       new_component_0_write_to.conduit
			reset_reset_n                          => avlm_avls_1x1_inst_reset_bfm_reset_reset                             --                          reset.reset_n
		);

	avlm_avls_1x1_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => avlm_avls_1x1_inst_clk_bfm_clk_clk  -- clk.clk
		);

	avlm_avls_1x1_inst_new_component_0_data_in_bfm : component altera_conduit_bfm
		port map (
			sig_conduit => avlm_avls_1x1_inst_new_component_0_data_in_bfm_conduit_conduit  -- conduit.conduit
		);

	avlm_avls_1x1_inst_new_component_0_dbg_data_in_bfm : component altera_conduit_bfm_0002
		port map (
			clk         => avlm_avls_1x1_inst_clk_bfm_clk_clk,                     --     clk.clk
			sig_conduit => avlm_avls_1x1_inst_new_component_0_dbg_data_in_conduit, -- conduit.conduit
			reset       => '0'                                                     -- (terminated)
		);

	avlm_avls_1x1_inst_new_component_0_dbg_input_en_bfm : component altera_conduit_bfm_0003
		port map (
			clk            => avlm_avls_1x1_inst_clk_bfm_clk_clk,                      --     clk.clk
			sig_conduit(0) => avlm_avls_1x1_inst_new_component_0_dbg_input_en_conduit, -- conduit.conduit
			reset          => '0'                                                      -- (terminated)
		);

	avlm_avls_1x1_inst_new_component_0_dbg_output_en_bfm : component altera_conduit_bfm_0003
		port map (
			clk            => avlm_avls_1x1_inst_clk_bfm_clk_clk,                       --     clk.clk
			sig_conduit(0) => avlm_avls_1x1_inst_new_component_0_dbg_output_en_conduit, -- conduit.conduit
			reset          => '0'                                                       -- (terminated)
		);

	avlm_avls_1x1_inst_new_component_0_dbg_write_data_bfm : component altera_conduit_bfm_0002
		port map (
			clk         => avlm_avls_1x1_inst_clk_bfm_clk_clk,                        --     clk.clk
			sig_conduit => avlm_avls_1x1_inst_new_component_0_dbg_write_data_conduit, -- conduit.conduit
			reset       => '0'                                                        -- (terminated)
		);

	avlm_avls_1x1_inst_new_component_0_dbg_write_to_bfm : component altera_conduit_bfm_0004
		port map (
			clk         => avlm_avls_1x1_inst_clk_bfm_clk_clk,                      --     clk.clk
			sig_conduit => avlm_avls_1x1_inst_new_component_0_dbg_write_to_conduit, -- conduit.conduit
			reset       => '0'                                                      -- (terminated)
		);

	avlm_avls_1x1_inst_new_component_0_input_en_bfm : component altera_conduit_bfm_0005
		port map (
			clk         => avlm_avls_1x1_inst_clk_bfm_clk_clk,                              --     clk.clk
			sig_conduit => avlm_avls_1x1_inst_new_component_0_input_en_bfm_conduit_conduit, -- conduit.conduit
			reset       => '0'                                                              -- (terminated)
		);

	avlm_avls_1x1_inst_new_component_0_output_en_bfm : component altera_conduit_bfm_0005
		port map (
			clk         => avlm_avls_1x1_inst_clk_bfm_clk_clk,                               --     clk.clk
			sig_conduit => avlm_avls_1x1_inst_new_component_0_output_en_bfm_conduit_conduit, -- conduit.conduit
			reset       => '0'                                                               -- (terminated)
		);

	avlm_avls_1x1_inst_new_component_0_write_to_bfm : component altera_conduit_bfm_0006
		port map (
			clk         => avlm_avls_1x1_inst_clk_bfm_clk_clk,                              --     clk.clk
			sig_conduit => avlm_avls_1x1_inst_new_component_0_write_to_bfm_conduit_conduit, -- conduit.conduit
			reset       => '0'                                                              -- (terminated)
		);

	avlm_avls_1x1_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => avlm_avls_1x1_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => avlm_avls_1x1_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of avlm_avls_1x1_tb
