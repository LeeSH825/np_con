-- test_tb.vhd

-- Generated using ACDS version 21.1 842

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity test_tb is
end entity test_tb;

architecture rtl of test_tb is
	component test is
		port (
			addr_master_0_data_in_condiut        : in  std_logic_vector(7 downto 0) := (others => 'X'); -- condiut
			addr_master_0_dbg_data_in_conduit    : out std_logic_vector(7 downto 0);                    -- conduit
			addr_master_0_dbg_input_en_conduit   : out std_logic;                                       -- conduit
			addr_master_0_dbg_output_en_conduit  : out std_logic;                                       -- conduit
			addr_master_0_dbg_write_data_conduit : out std_logic_vector(7 downto 0);                    -- conduit
			addr_master_0_dbg_write_to_conduit   : out std_logic_vector(2 downto 0);                    -- conduit
			addr_master_0_input_en_conduit       : in  std_logic                    := 'X';             -- conduit
			addr_master_0_output_en_conduit      : in  std_logic                    := 'X';             -- conduit
			addr_master_0_write_to_conduit       : in  std_logic_vector(2 downto 0) := (others => 'X'); -- conduit
			clk_clk                              : in  std_logic                    := 'X';             -- clk
			reset_reset_n                        : in  std_logic                    := 'X'              -- reset_n
		);
	end component test;

	component altera_conduit_bfm is
		port (
			clk         : in  std_logic                    := 'X'; -- clk
			sig_condiut : out std_logic_vector(7 downto 0);        -- condiut
			reset       : in  std_logic                    := 'X'  -- reset
		);
	end component altera_conduit_bfm;

	component altera_conduit_bfm_0002 is
		port (
			clk         : in std_logic                    := 'X';             -- clk
			sig_conduit : in std_logic_vector(7 downto 0) := (others => 'X'); -- conduit
			reset       : in std_logic                    := 'X'              -- reset
		);
	end component altera_conduit_bfm_0002;

	component altera_conduit_bfm_0003 is
		port (
			clk         : in std_logic                    := 'X';             -- clk
			sig_conduit : in std_logic_vector(0 downto 0) := (others => 'X'); -- conduit
			reset       : in std_logic                    := 'X'              -- reset
		);
	end component altera_conduit_bfm_0003;

	component altera_conduit_bfm_0004 is
		port (
			clk         : in std_logic                    := 'X';             -- clk
			sig_conduit : in std_logic_vector(2 downto 0) := (others => 'X'); -- conduit
			reset       : in std_logic                    := 'X'              -- reset
		);
	end component altera_conduit_bfm_0004;

	component altera_conduit_bfm_0005 is
		port (
			clk         : in  std_logic                    := 'X'; -- clk
			sig_conduit : out std_logic_vector(0 downto 0);        -- conduit
			reset       : in  std_logic                    := 'X'  -- reset
		);
	end component altera_conduit_bfm_0005;

	component altera_conduit_bfm_0006 is
		port (
			clk         : in  std_logic                    := 'X'; -- clk
			sig_conduit : out std_logic_vector(2 downto 0);        -- conduit
			reset       : in  std_logic                    := 'X'  -- reset
		);
	end component altera_conduit_bfm_0006;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal test_inst_clk_bfm_clk_clk                             : std_logic;                    -- test_inst_clk_bfm:clk -> [test_inst:clk_clk, test_inst_addr_master_0_data_in_bfm:clk, test_inst_addr_master_0_dbg_data_in_bfm:clk, test_inst_addr_master_0_dbg_input_en_bfm:clk, test_inst_addr_master_0_dbg_output_en_bfm:clk, test_inst_addr_master_0_dbg_write_data_bfm:clk, test_inst_addr_master_0_dbg_write_to_bfm:clk, test_inst_addr_master_0_input_en_bfm:clk, test_inst_addr_master_0_output_en_bfm:clk, test_inst_addr_master_0_write_to_bfm:clk, test_inst_reset_bfm:clk]
	signal test_inst_addr_master_0_data_in_bfm_conduit_condiut   : std_logic_vector(7 downto 0); -- test_inst_addr_master_0_data_in_bfm:sig_condiut -> test_inst:addr_master_0_data_in_condiut
	signal test_inst_addr_master_0_dbg_data_in_conduit           : std_logic_vector(7 downto 0); -- test_inst:addr_master_0_dbg_data_in_conduit -> test_inst_addr_master_0_dbg_data_in_bfm:sig_conduit
	signal test_inst_addr_master_0_dbg_input_en_conduit          : std_logic;                    -- test_inst:addr_master_0_dbg_input_en_conduit -> test_inst_addr_master_0_dbg_input_en_bfm:sig_conduit
	signal test_inst_addr_master_0_dbg_output_en_conduit         : std_logic;                    -- test_inst:addr_master_0_dbg_output_en_conduit -> test_inst_addr_master_0_dbg_output_en_bfm:sig_conduit
	signal test_inst_addr_master_0_dbg_write_data_conduit        : std_logic_vector(7 downto 0); -- test_inst:addr_master_0_dbg_write_data_conduit -> test_inst_addr_master_0_dbg_write_data_bfm:sig_conduit
	signal test_inst_addr_master_0_dbg_write_to_conduit          : std_logic_vector(2 downto 0); -- test_inst:addr_master_0_dbg_write_to_conduit -> test_inst_addr_master_0_dbg_write_to_bfm:sig_conduit
	signal test_inst_addr_master_0_input_en_bfm_conduit_conduit  : std_logic_vector(0 downto 0); -- test_inst_addr_master_0_input_en_bfm:sig_conduit -> test_inst:addr_master_0_input_en_conduit
	signal test_inst_addr_master_0_output_en_bfm_conduit_conduit : std_logic_vector(0 downto 0); -- test_inst_addr_master_0_output_en_bfm:sig_conduit -> test_inst:addr_master_0_output_en_conduit
	signal test_inst_addr_master_0_write_to_bfm_conduit_conduit  : std_logic_vector(2 downto 0); -- test_inst_addr_master_0_write_to_bfm:sig_conduit -> test_inst:addr_master_0_write_to_conduit
	signal test_inst_reset_bfm_reset_reset                       : std_logic;                    -- test_inst_reset_bfm:reset -> test_inst:reset_reset_n

begin

	test_inst : component test
		port map (
			addr_master_0_data_in_condiut        => test_inst_addr_master_0_data_in_bfm_conduit_condiut,      --        addr_master_0_data_in.condiut
			addr_master_0_dbg_data_in_conduit    => test_inst_addr_master_0_dbg_data_in_conduit,              --    addr_master_0_dbg_data_in.conduit
			addr_master_0_dbg_input_en_conduit   => test_inst_addr_master_0_dbg_input_en_conduit,             --   addr_master_0_dbg_input_en.conduit
			addr_master_0_dbg_output_en_conduit  => test_inst_addr_master_0_dbg_output_en_conduit,            --  addr_master_0_dbg_output_en.conduit
			addr_master_0_dbg_write_data_conduit => test_inst_addr_master_0_dbg_write_data_conduit,           -- addr_master_0_dbg_write_data.conduit
			addr_master_0_dbg_write_to_conduit   => test_inst_addr_master_0_dbg_write_to_conduit,             --   addr_master_0_dbg_write_to.conduit
			addr_master_0_input_en_conduit       => test_inst_addr_master_0_input_en_bfm_conduit_conduit(0),  --       addr_master_0_input_en.conduit
			addr_master_0_output_en_conduit      => test_inst_addr_master_0_output_en_bfm_conduit_conduit(0), --      addr_master_0_output_en.conduit
			addr_master_0_write_to_conduit       => test_inst_addr_master_0_write_to_bfm_conduit_conduit,     --       addr_master_0_write_to.conduit
			clk_clk                              => test_inst_clk_bfm_clk_clk,                                --                          clk.clk
			reset_reset_n                        => test_inst_reset_bfm_reset_reset                           --                        reset.reset_n
		);

	test_inst_addr_master_0_data_in_bfm : component altera_conduit_bfm
		port map (
			clk         => test_inst_clk_bfm_clk_clk,                           --     clk.clk
			sig_condiut => test_inst_addr_master_0_data_in_bfm_conduit_condiut, -- conduit.condiut
			reset       => '0'                                                  -- (terminated)
		);

	test_inst_addr_master_0_dbg_data_in_bfm : component altera_conduit_bfm_0002
		port map (
			clk         => test_inst_clk_bfm_clk_clk,                   --     clk.clk
			sig_conduit => test_inst_addr_master_0_dbg_data_in_conduit, -- conduit.conduit
			reset       => '0'                                          -- (terminated)
		);

	test_inst_addr_master_0_dbg_input_en_bfm : component altera_conduit_bfm_0003
		port map (
			clk            => test_inst_clk_bfm_clk_clk,                    --     clk.clk
			sig_conduit(0) => test_inst_addr_master_0_dbg_input_en_conduit, -- conduit.conduit
			reset          => '0'                                           -- (terminated)
		);

	test_inst_addr_master_0_dbg_output_en_bfm : component altera_conduit_bfm_0003
		port map (
			clk            => test_inst_clk_bfm_clk_clk,                     --     clk.clk
			sig_conduit(0) => test_inst_addr_master_0_dbg_output_en_conduit, -- conduit.conduit
			reset          => '0'                                            -- (terminated)
		);

	test_inst_addr_master_0_dbg_write_data_bfm : component altera_conduit_bfm_0002
		port map (
			clk         => test_inst_clk_bfm_clk_clk,                      --     clk.clk
			sig_conduit => test_inst_addr_master_0_dbg_write_data_conduit, -- conduit.conduit
			reset       => '0'                                             -- (terminated)
		);

	test_inst_addr_master_0_dbg_write_to_bfm : component altera_conduit_bfm_0004
		port map (
			clk         => test_inst_clk_bfm_clk_clk,                    --     clk.clk
			sig_conduit => test_inst_addr_master_0_dbg_write_to_conduit, -- conduit.conduit
			reset       => '0'                                           -- (terminated)
		);

	test_inst_addr_master_0_input_en_bfm : component altera_conduit_bfm_0005
		port map (
			clk         => test_inst_clk_bfm_clk_clk,                            --     clk.clk
			sig_conduit => test_inst_addr_master_0_input_en_bfm_conduit_conduit, -- conduit.conduit
			reset       => '0'                                                   -- (terminated)
		);

	test_inst_addr_master_0_output_en_bfm : component altera_conduit_bfm_0005
		port map (
			clk         => test_inst_clk_bfm_clk_clk,                             --     clk.clk
			sig_conduit => test_inst_addr_master_0_output_en_bfm_conduit_conduit, -- conduit.conduit
			reset       => '0'                                                    -- (terminated)
		);

	test_inst_addr_master_0_write_to_bfm : component altera_conduit_bfm_0006
		port map (
			clk         => test_inst_clk_bfm_clk_clk,                            --     clk.clk
			sig_conduit => test_inst_addr_master_0_write_to_bfm_conduit_conduit, -- conduit.conduit
			reset       => '0'                                                   -- (terminated)
		);

	test_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => test_inst_clk_bfm_clk_clk  -- clk.clk
		);

	test_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => test_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => test_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of test_tb
