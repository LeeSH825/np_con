`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BZuLUnRBD+r57HjzrB8/gKYCureh12IvOjK3U87pgMUZUum5BKk9ZYkuwOEd6AAA
s3E5Mp1swNMz7uCaPPKcJwiivz8UOI6FFob15LZpSMhT70ZIY+k5cDxSf7VWHYu0
jUbvVWvO7PzTsU7s1SN5LT+iE8Z+6cP86iie3/s+JqU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 82944)
r0n7RdhJS58h7FEYQYi9InYv2wPJpQbBpHG37VhyglI8lNqHaU+fmkLhE2AyeoXB
ntbv7aN2foKf4mGLOPXjEzxDOUm5EfTEe2X2YXaZ10y6RSwK19+s223T8R5CWCRc
hu2EXhWb75q6NCz1NZpStvK8g7A/jaJHudoPY438V1NSwFc7wBQkeNzD1P3fqtgf
2/rojlVpXknpPPTcpPZiLHKFlS1DNQ4Eq7G8OaBC3CTaQdDFILVD2d6c1ULCWT7d
qlxPRSOL4p3soFhRAO8zUWOcEPyoQr78NtoZRKLSv5+FhWpSMHWDOYdu+VzXq459
cfeKjXOO/nVeCkNzP8Wu4lqZal/SenlpyRtlnMpBihrrbbfmcdRbXmoDH6kTuIFq
jXZMyrwOsOEqNx0U2oMmv6xPak+UjI9r0e3HYWA0vGJGyY+I9k8BgC2LFNb0Agji
qBt4Rdt7+yCEKMGu/MkkD/u50Kx+8eJ3t0TaSYVVwBHNgZMGHrUNY0rGjS4dfbqC
rgBTgyaar1eVOEj7LqfrQA6K5scFM0FCEMMVjiM2kvOmUiDBJfC26AtsSSOUekGp
8+Ti4bQbYoCxRSvmSefH3iR9M+scoslaUnx/mBn7pSWSGLk1LSgJiWTo1Vn1QyTy
cgDfwL4MwMZUaiziAb9Kc+hOVa1FKaxUm01s3VNL/oTTuDSLGYCANic8ztxaWP42
LOtXtqzUf+1JuXEdv8J7lsO1mYjx/ESIH2Qt9zNOtZ8OraAhdiTJ37JyFHCjKTaN
8ZpOwDF9yCdVV9im+zT3/kRsSZv4vC3l1nbl3Hun+bu58WD1UPbP/7PkZMDUEue8
RxiFgdkZQu4YAZ2eI1coGg1FgOD1ytHCHg2y3os25WE1WnRHS3gOJ4RnWt/QTubQ
KWfRN4NZHWOfv3WouXvpDKvEU+dx1Q37ZbNwWfBamWZAuHmvYSiEyIbt1Of++mRf
yPkNf4/I2bYLJt0+vZ5pNDAsScjvIZCgz7klAiQ/QXCVE0hIqGktHd8ETOlQxly0
+/uS5xtjIEOALHN04xM7AONpH69xMsbJB9kWHhC9Qytf8saiBj019MaxkeBHxynM
ERF/rUzKrxlKlt6+vPoFtoo5YOPGbQxOFbrHb1SCr2zbVz6S9JasmLeJ1JAVHy4z
rPboV3EhSGSLYcStpX+t0Yn9VOxFF8rjqx9jmCovc8GinvsCYiyGJMLajUWiTwJS
kp/3zfD4oxPS3ffgoDmZSJdsJd3dIxIr8iW4vlake3Y8xlb3nqMva3C7f2uXvKWV
9fRt4CNAwrieklUi6B9s4iY4r3qhHwcsAxgb88Na7tyRFoT+zOayzY/lGX6iX2Ap
nM9p1Btg/LudUjkCBe7mBMmepJsYUrDbKbmkGTcrakH6ieETrf4/pYH1mJiSQxTS
CsqeUS9n8Z/ZI/dvABVd4CPltKvv5g51TMjJjGhEUwwzTEgn8A76xU7YdDcsfNjP
blE3kFeLs3NNab8ttq7zDYXkjJE0MGrOiE0cOCzAZwCA6/oUp9z/GhKvNRHw/DL7
56OQHdYNyz/6k8YXfj2iqBhdOp2jDq/QmnaMhfVCSnoYg21W+XJZIO4dyaYVRL2B
lY2khjJGiCprREag3QM+pGULZdfIc7Rc8qlQr0Ht7CyrQwX+i1Gv63fnn4ao4F2Q
9hpWisKpzDxKTjvKxsfRK/NWL6CxtWtWO/HSMH7N5MVCqLSQreLXGuORQO7bRP/O
5GMjIL1iWSgghpJTFbCovyxwn9SVyyilZ5r2IPdQSbDSuQ7BQooh/Q9uwIYcDf2B
BpnlhvGM30S3nyyPo/huMgrjYk2ksZ07n+CoXjWN6RjP4RbxZbCHdZYdTzRDHCRJ
IBT6VPeKWiRJZrGFiusg9GyiIGYdlneZT9Pqyytl+JYA4G6MQFwM/MSFfaRzd3b5
gtRkDkZ0BVIhFSMqRYeLaGU6v9SCDfxWRny84Wyu47YXYSV3ZPXXxcr7iaZbgdRP
SjTcz/92jlsMwGvRtimHHfoUfzwteBKUKLAxXHsfXVsQXmggQ4w4wjF3tj1YuOA7
IDGAykq6KA6zAEEYVQ3CrIyJm1gV7ty6SmeN0lqXi3hqga1fIokT3n7QfePa6Rgf
v9t8/9xQiCTxU/EexzhVwh00d9xCPSOhtBEVT8nWP3KdXQzwX2FyDOo3+EQJVQcE
4LT7maLtQfIblpjZloWvy2by9Xc6Jdu0FNPXRQnIY4eUxcaJ18a5hO1UwD/AwZTg
jneHsQfxobExc/iYqs07Xz3xUQV1UEqxJlGnCHsaKjIThBYGVyGAeZZpvgkO9V+Y
bIyFhuTrR9vzf1szJvujxUZgYNabMj7KnoL9fqGpBIY8dAlOKSpLQAchOnPGcCg+
9RJ4X6W6pb0eEemRw8pu+b9EobClmyUgrcNhxLjGH1E3nU1lBQk6MmWGFcDnjQJj
nbZpnfhcERWhCKCDW9Ks9LTeRzlpVACDlrmqAgZs2XGifkhJcZkf0qTSQV3GH4b3
GijRJZU8YU6FVWftn57fid19Fi9P6miox7Mv2NMPt7GlcxQmOzWfHam0KJJpUNZr
orKIkFZSksgbMb+d1G76yBvKFQsUDS3PLSHEvvYF2imayZ/yWR9l0YqDZ9nricen
6Tq5xrq1V338eXJpag4QlEja8ixy7hogdr9ZSkSX1JXUHt2h+yDT0iqtKVvkAbNq
Qei3ok+2qN2GfDtuWCeXsJiN8uoGCsgDfkV12MWjXjxg4JlKK1m1aqhzTelmeONT
0qiSw/frYUDOGRSusLcOG42HLcotvYra3C1aAFfEHPvalAqInGzEUFjQXLYP+nWZ
C57f9g6UEwwP9c63bzXrjpMsE32oRWmpQl0HFImEWLaoBcFK9E6o0g+n8vLuI65W
03VSmRQc9WJwHjaifLsezFPJ/0SgS2z4rUmp8fNRizHS0BDQEJdxnOflB//wn22y
0vc5rLv9pGry7zpxEPmsh+7OVc0Rro2KnjKm0qEfpwhSrO+1CUB/FCCzlk/T+LHv
bEeSWfLrvMGmfu59fFgZIB5wgqxuwTwwytrgB+FfQmybQV/5w9+RjN+n0p9Se7gA
7lagMeIlJeWmaM7YU4fG5GqQEegGbb3AtCa76p2Y7QWAJCl4/TMG0z8ubyUssGrQ
v4aZLp4R5vfXfJdlg5WJXuLrsQQlw0IWTVn05wVrFXFQ6bjw3uX4hnraVwlC5tBB
dDl+ibZjyZK1d9VWB1xYKTzbHHVA2IeitwIMEM2bimNG1Dj635QpzoOkmgCnc0gv
lTL6sLfEkL5vWXEokVymYL8SgzSsM72m+PMKgGSOLkHgSr5Yd4jFGx1IMUK32szE
fC3+tvZ8powfvnfZ42bUgF0cA/g9kMW6nvAhjp7Z43EjsUzhEWpz3Hw8ANire1cn
6Qn7W9uYkTyYoswsVwMFcEW7PpLjVVcRebN8ZSwHVlIbqJcfJQ16V5Xk6uNJW5yx
LCVXmkXI83I0mq0tONyYEJi+6hiU7VykPE1ETch6qTobB/Zm2PC7H9zo2qFN+8Qz
pltBNUdoLU+7nXjslZcy/69+QcGvQ7Kb3guQ000OIjZs+SNeOEUOvJD1fj/iMUQP
YcYr1J/zOP/vAb+AvfjBFFRkWS3lG7+srjFBMpbGhsPGf2vGqLtNSkdyS5nILH5p
RNuETnPvcDndz8EuEWZ0F12YTriWdmduVcGIxserEZduLVUGSsRnKoeIheCAo59c
Dk54B3MW7SOGB7GJjYEKt9CBCd1o9ugrnCyUzkJufs9JaHOewbAqSQGitbYeVu3k
40Dtm5yo+c9E5Q4lvt6yOxAl29/ccIOXWgS9Qu2nuq9HgoU3+cFk2MxoTMp6UDys
PF7aVLaf1SOa61IZSCS2Nb8y8cEhqUPmeW3hKj6KIjyeTjqU1T6xDq/JI/r6Klqz
aZyMiPitUVce62CYwafxvixEUWuyGh4cUAsct20AcIRev4IihcRRtfDswnS3iAVR
a0zh+WZEHs1B9c9bJVn8jXmJRxhU4yTNgCaVzHA2NnogKdWiy/0F9s2rOPj1fIYx
eOjf9Y5nfim9oG65ERR/5iUa4LtT8saVV37EiXYwP6xuBTH7li9rzvdMsH80TiEH
+DM9tSRzyZ38Q4b2PMKRWeLgYNSpbT5YxOlq2tuE3SEsCy5gYcwmn9PusKqTHFha
DHU5njfNCdC4veCJs7qMqlHcNp1FX6q19VRLbcS1WwvcdR1ZaqYWhs/NmA+SjSam
P5UehaKCUaqhq1rpQNReg/zQHVL1xlfV0gnsChhZQt1ZFMODREyJFnkguTUwUNRb
FFI8NRdbJiDJFiya16AsVF5sx5pnWbjhoD0S9esQcUSSPpSnDKwnyExQAfoH4+aP
tAsFBfXPiTPJ/okPaiYHG49sBK2hknnbvflGRizLXfsgWiZ1Azo5n/p/IKSzE2I1
PoSu+YW53vsJG8co7Y9qw/56P5+rjrzsiKOIGzRlk52WNBB2fJ/onkdoQWNOB8ac
3nlwCQr7jngU+N11dMYBRcCrSKnApJTubcGl6tZUtMPqoxamGZGAMJJA5IBm2xfm
yCQEJwAOx9pJB+FpZOme0S+qlDcntrgCmIWbLyov+ugE8OdL7azxjSfungFT2x+T
idcp+oOKbYnlTqYaxZYggZcxvoQP3VUIR9B/zrQrxT5nbcAf94RZXL2S3spgReLq
AhU9dCYBm9jC0alGzgQAyY1qVzhJVG8gGs2Vs5GRdh6nF2cnT9BS6N4sQEKIjz95
EoEkNq6VHeX3rCIOyqaJMoIZEHeSxHEFN5wnGXokA5TCqgyjp9n1Ly1+ETIyS/e8
Qb5nxGFnoVWTrMXimFtCgcYeDqf60aWJOlUgBcfTjIEi27ttEE+BnjTR3YqWOod8
zrqn47V2C/5tcuUjFiPl0E26OLtlLCPDKbdt+j6FqefwleLQFe6kdgb+FCXd9mp6
ZGH2qrsmcDM7UiDceFU3BsUdAbAOJYYz4jkmFHutJ8kESrhvxF6Gkl7WjreKf0CY
sVpxyZLKUAPso92nWuKCeTAVq8kLmG3a5qOm4QLNAaXqLaamiZDSLxXTO8PuaCG+
eSLpbEZ3NhKvoRaGYRz/YGETVuc1kLU+bcE4JBCTe9dhT+L6UijnS9a+gpe+YXcA
Om3H666fdSlwbVJ1P6gaxLTd9Zi7bLBW6Ew/BaI/G5Jz/vAuIQSwIwMw945fCwFZ
x73RKbd4wZXpFR//QzceS6O9M8f4WLMD7PJhAlVFhRWiBR2bdtQcpJnsltanbnBx
wNQYRZzG33AU37WQyffMPmwjNTnqYh/7GlIvfBWmFeM/rZimb2/hu5ZtjUYWvpwx
tXlsnE6JngUClzpsRX8SrVDEyTIdhkb3NdpBjgaOVKyqn3mzxOKVXtgY6ANDQOMM
uiQT4//kC8o1BxwMj2tPeuMFWR2aYRTewgN+Hq89SHyI0HR/t7CC2gk7XUSq3YEX
1vonCYG0GxpPPr4WRpBqfUtk77wyXsgf5k+efpEM9HzP+0diQ5qtKC2mvQ0SUzKS
O/4XInKpqMyzaMnYAk1eVs89UY0Pvum9mdrnM5dv1nYg+wKkhlsJ7SH2l3ztRix0
njamQ3kj6ed/L4USOlZZ+BTAQOBy5+9691E+ziJHAhuyt/wS6ERg1rVijBQ9Z69C
sew0e0BteZkLSS98iRMspm640Ek+jvDyqSUBe1URyZsl2dhkl3xupEOsHyPmeXLA
sKG3k0OG24zysoI1AmjptoFulA09Bv1ERnkQoj4Xa++nxNoHiqwCvkS+yDXuNlmd
nJzWEwUIPkx3W7Ro8pHVfRayZIiWZX8CdvVi+0vRV06ZYItKHl4E1TRvVkqqAlij
BPb5geFxC3bIrYGNiq5iqqo/ck08+fBLNu+HsUjMZs4JssMG/8Cg1gcXwufrPePp
jq76ts/JeQKpcTyNtZVAtRbzSBYliu9YQaXtfOuh2r2KPT4f3catciBgY0uEDjdA
0Yplh9rpjMNHIYQAbFJnPjh7QzvZpCR59djnRw1TMqB/a37QZdPkNC9LsqDP5MYv
TCrrFB3ZlHkCavylPifJZiIwFrF8vK9I7jgfvVwLIgbFNlQwfZHZDitc9Gnw3ug/
ROY2n/mqJDuhUIEVRChFj7W7SN7d1IHRrHm0IkjOVycjGLtcsWhLmwTcPtueazJt
oTYEsCefelEJtYC3LRsY1WmIAoNB7KgNCwcLV+FEdx5Cc2ThwRn7S9xllYnzTZmA
kHDBUpPfSOPaNwIRvifEW96CRcQA4SAaa59ssd8vAYgAjshPOOsTJttEsdNCnFdv
qT2QuSRUj5Nnu9Daeh5ZFgl7aREw8PAPB8geWi+zHx7ZWzKu5TTQUjU2q/N+Df7n
1yMbrg/T2g97VAhsoziWJ+FBO3T1hi7nK8NdRHafFseTqDs0qOXnq45W8YFFR1O0
A2k1P5gu03Xlz0Tl+A9teXY00mid6G+8l1Se9f70VwYO3MIz9jHN9RidIobH1W6z
2IjrM5a7XBNHdNVUozm2Srkpi/fI/KvmPslV3LvB5jXPBDDaDeEUIGtQksnCNEjo
73EI6B4IyrV4QwH7rOVDl/zLmxHXF/IE9mC3cuTrjY90A7F4JESeHdunCHO4hWFC
KEbzKh5Rk4sWhJX4ahbFaBKzpp0wGO673+RO3qJZXow0cVG98UQrQ0/EShYyvAjb
atOky9ElnsIFwj0YwJ6nOFlYF0/esDj0KLlMQlBiaYiJ5CPzHerNpCluOXzEqY++
lY1N0HOoY0BAa1TKWrKWTw9FfEIktw0l0mWrLqzZB21vsZlYRN/6GwcYynI3NRsw
x0MF0HX0qHRsG5uPz3P6c98WnmLHq/EJYEi8UP56GtFhCMm4pJCgWloVf5nyf7Dk
paySzooRFHuTHpz7MBzXrrzG+WZzUeo2gM7U1tXy8c7eqUlIfNCJDaTvd/xn6++h
yaCXd231aqdO5+Za264FdbIIwy7irxdYb8QD2wazXP2wvKrCEhIJPuihdsH2KKHT
+i5rWt+s0K6LAuzc3GCfYqaWIIXrheADBaQZ7KLc3nPw0+CuEzqpJxZ8AibA1jXV
un+CEXdm11dyn6BFz0S41W6fpibqTZ2yzodpmhs8zfpuCKQC55Y1b+guC++yHMvJ
HF9Li2Dy4ur2znBsR4Ugi9tpPc80KjnBLORYvt4axuWBFsVh7EQTHs/ZGMC6mVQ8
zNfZPUjZ9LsgN7lHpkFaIpfVQX/nHTQnGepr76FAdhyvnh5AdygFO07wQA7EZbgy
l/v6zI7NPclthkSozmpiF+/xwCWYVvq7KiPu6cjORKRBKlnfQe4IpIj3dduf4Wbe
wof9p/3VI8l+0+tB9Z/5jmL+8L4cAL/50VXNWi3ZzAC3Dw7Z/cb2YRgsiRdhJgHz
0byriiNhIANIuV+0kIn0NrWSVjuNRAk/ax2jtrh9FGgiJmSVL20CyAolzkec0GdR
NZhphEw9t7BpizBZ8ZHsz7FhOO6uSCgWQlF2OxdH8Tlp2uDzcycdyA0o4q7VPPpk
866U7LmnKmtRvglCJ4FxYBMgJA7jPjesO0fT1QHtovvVLJyNRe1Qh4QM+7uX0fpv
qNMXDDpqQ8uBGb44/8auEHG+dMu6Aqx1X5tOom9TFWFWLZvk68ym5+HiE/ojdA64
IR8X19iBidKKFbr1i+pnFbZsgWhzZSqUL1K3X/0yATEu8Fn94Kn/+/gSArnE2xBl
mGxnBukFjrqa/ZZcrB1/junDG9KoHrrL0NLiwmDX3c6YxzKjEVn3UfglgQ9eQCiw
auENqCgLrGnkC7LmYXv9zcC1GUKGxNPffZ6HxQTcSgd2iBdHg58/rFVEa91x25wR
MqAPYEWJgH/iIVsqS46nxMfMp9yS5B7vrKiH/xj/nWJlKpw458Xa8NBfxJ2dAxBX
Y8Wkq5eTHB6S1+0F2CdvoMnysCsQaZ9hB+LfyeG/1LK4Y7w7XFoSqVRHYQXC5Nto
iCARtb1MWx/Gwz+9823RO/0WUW89PABl7+ZaGkDyZy5hKEbqcYAIJPVuuJ2DkrVr
vFnNUTNPQs/meD9A9C5DpuabCDWjpGmnN96tlRyDMxPWUlejapOvRbGdfXSqgklT
uX+fxboDdnaYcSK5Ru/uWoyC7GTdLY9+7+UsvniV+ZssDfUrzhY+anLpP8UIuxiL
sEWBHw6wxpKfauRIpUoN2fPYBicnDEV+xWrvQ4zjT7+iLFxujpiUHM37NbwlabGL
QW/GkLN+/OpeVJW92SIjO2uMaxP+P4zcQsz2+MKvIW99s7ZOsNEE/dOztuatTacm
Uyu8gHNuv+gd9OAzHME+nnydOZjdAmcDO7+EqI0s1BOuPGjHkc8SJaQ/y5Xxc9yT
aZLaC2n6ckgCF5I4BnQZDD5oG4xSg9g57OVr027NAFun1L0At6DSNgTslttRYhnb
WAhaASQVIgeL0kL76tSZYlromfWp/fsMcLQvodxUg8ntM+QxugPHK4l+6L8j/uO4
auuvbNv2EOjpIsbNsGW53mPFWqIyN7smxzFU5jdhQDGfQ5xBoB0zNaai763HQP7V
H6xHRUWjPOPU3ewUn74xrw70xWN+d1TNoAthvWhiMc1c9o8ZULx/0SP40Um/j3M8
GA8h1S1Zxn7C6uB/7h/dC0QkIElRAkygwpVuvwJqzS597XHS96+O6TT5qJ7FOnNr
RSazyAviQiKlxK+I1dz7DzNtjlosupNcvPpuBW/IrnuNuGyi/Fg9RESmepCsgoEV
rlGXZ/3lmc1e9SGLjyXE5doeZb64Awa/jMcLJYRSuJjOarqTyz1nLcWVfWwfMveI
oGCERhDTne54OZr7MOvUmm7Nza2RhMv0T3XZLyFfD1b/HptScK1oZTwK6GOh+DvW
RzjEv1LEaLrb9NSCb809UAvo4PeHvxLatvPAGgH9QPdBvk3q+yQxcy9JcU8gb2Tu
BMB9w1s5qvofrtLLnuXOyOQhCP8mQcA5R7zg5ansvL4APurawAFK5dNmizZYDq20
x9Yhi+W5ETLIwDBxUo8wczhdCaX+s2ZEyNXRm66u6B4WBFHkdDugtqtsQ5mYCHtm
y7m0NHJdokueXZbjz1rrMOGahv9K8A1+Bhl1C6Ci327D6dMLduApZOlAocr3kupQ
jmwKwHWnKMvG25WxwRCyLErDvlxrvRnAXjmNTO6fx7xA7tqqcsHjojugaBGQcfjK
YBYq37QKHQfT3hOe962bswGA1ecItdhgZkINTr8cFER+yblEMVhXoUC7iXS2VAye
2zxgaWC8H2eI/Jqbwet3PHe/DxNxi613O5pSL4InqZ8VzefcBgZnlC10PzxR4v4C
Q6VIX0On54GFgxK5G/BEXrW1FkG0V5oawjmXQXPDVw0goyj5LW4PYJktJ+g4rgRq
MHODq7O/jy4Sh/5pAg8xuMGUCZUY2WWazVUdofVaWgso0gsk2wIig+plP1Vbt6AQ
TKC4bIqi63SYGONs8HmtGL2M+p77wvZPk9Egv1n07fBwZqyrcoz0zPPDJPBYca9M
8pymeEzbJQd5ryifLRrvJaaYJ8vDzG7jWqmw3P2rkChaq6A5dobsr0WpfUbdw/ER
ILyCVKit+0Kc8N9UbsJxaMNNMl9qOgtcKd1vg0KJ3Nw6iiXrXQHgf4ZeuqWpiJOW
K4xvkbcwHD4uBEg9dRkO811vTQFq5asEYJb8gzSR3mJRQ/uB0ORVr9xbNKYTFLfD
oYFTU297AuFDL8TgRJhDUavCOCkLb7z93PKmyI6ptl4IKbFcWzzZSZGylyLKaGoK
a/MbY3UxM+pTssu02+QCquSw21FYh5gCaG9YHvunmQmJYZ6i3S1hlAa7zO/7JuS2
rTuY223h/x5b+yesmoWLI4JZjkAwigZMjaRIOY6Ml+2nZBb8/ebHnxw+H2bIkhJu
LA9OLcnrNdFZCAD9n2EhbTi4pR1p/X2Q9qOHv4S4EeX451ZdlNlbK48zZ7ij9E6I
oRuh1TWrE1DZYKFl6UzlztpnyYUAAHlnRi5jDZsHf5qpyvXAeYSUbcwBL1fIihp+
CpXFJLDVDV23V0KnvEdQGBSw4FY3IUQBJDTqhkjrBzqfra+pT6KUYvxI1o2/iZsF
aYhAHg7p8Dg694JIC6/yL2PxIozvPNf1J9XwVc81/K9IkQ28I7w9dfMMXMtY6R89
wZHRy71GCiNFBb3oRI0/FuJdz3JzPuyOgE5f+/fDPYpSUoE+50GpmODISGNjEmCy
r0i5F6o7K+cpUBz/JdNYZq4Smq01N9IDDyS/IgnV2UF7vyGJ+uCin6wWczDhmBJP
REoXYu+MhQm1HuYcbVOBcMAKUCSe9/GOyGCcO8zqz+e14J39x/eOXOiAMiV1EukO
1cF4qt90VOQF92xBAN6Ammz+acp7dT2aKJxJR4LkWJJrigz0SBAsB9gl90WBjCKn
/jb2Esg+T1pY/NefDChcFAW/IapUANDcxNgBjGkdZIZfuAcWtr50+thsW2BtUw/c
a0atvRCafkXWbWzrdUpU608HKyZh/OymSeUkjLSzFZxM9B31Oc5KjKysEsQC3oxi
396TfKVX8sLFFv2GRQqmYY75LKv3N3Gzv1Cnzf5XFttMTmxRLBPZghhcPnCzHoZJ
37S5CLpiFYoKZ4VrOOxBt9DcpVT8Wpx+OGfqg3X220O/vTVaL0aFtoRDpBnaHA5v
d/v1aFHhC17+0bKU5aSMmamx4bD8TufCom4N6m+ekM4ixYNC7bSeSpCfPgt2jxI2
axT2k0U/VWz+/XSa5pTFgdRZOeyGtGp3MXnm80HuYfHFf8V3O3ykqCSQB25cCJj1
lsjfejDYsfmaljL8U3XFw3nMPnJ96d+XwT6JnV4d0ed0zPekRUj6Co4eEQRE2sJD
En9xT61pneZSnruaZFYjpYyjbhVdtcsM2Au9Y4hMPkJ7J6cSQAzpAiexkN3IiIG5
XncIXaPEbbZ/SBc9R68OvJcjvETbV0egkZ7VrxvkrbwTNy7N0HIVgaeW+fJ0IAZY
jIp++azqcz31GagqoOZkYFEJEdSZpnwPvH9EGz7/BxAGFIocR1Cj8IDk0Eo5cuTT
3pzQogPE5Iu08ew7Zpn5z55AthVqfi+4ARx3ueQ4JHFlgNa24Na0NuFohZo33oqe
vOYE/LKtxo/1DY95IRZZCqNGNAtIG88u1p/jRtFZdvfzi9WLuAOsIQExD5s+Rydc
hc/uCcwtGQ8Z5/WvItyyNT3cspSdHoWkGlOKd7CLJOZ6l+HMgi8UREV2W/oH3/qU
qxIKh+shZatoudc2GPR0gJM7Pq2+3DiAjkECRcs7MQChcaVopldRiY4TBgXNSOMM
tnvTQZMngAQ3o9ZcPXt+3T6SovNVKPaDgEerw7MHE8iv/Gs0sUC7ozD5CrgTOmkB
9hDfXS2SxWKQtgspOJiBHBOCBtju2Xc/dW+GdRYdLMg8hF2Ge1xHz4AkFO9ouU2q
GcvGNhg+wtyVTm6LWVAbvx4/Iv71YGkzhVMFRMFX9AZfPClskHheYtpoQl7vYii7
DfipoSrd1dvZjhsb6eda/YD34jLX0CclOltx/AksQHwp65wsv5ckDGxNNRYLq4Z3
DqAMTnZOn7RUi3/nUHI/dK0t24EaSc5u4oWpQibsOSCeaezoAEePXFbl9FOX/gKN
j1fXBg3CqR8C/lvK2d028VS3a6rGJkhzxErHD73lIm2TzD2000B75qVlnhhQNgKI
tf7M/1z3zRYdAZkl5DKjr9OiBkn1OVIbnIUygjsFAhaYra1xgF4t145uEmUm/5dM
HxQtzLc9m1DDAEzAmZfalL0kyiHg261pWntJmLakBLLT/2H97suwvO3EHZ7SiyBo
qHN5V/LE7nS4qgYdDSHo1WNIFqCnTjVXYy3z+8gNqbsPF9fqePlz2Im0kGXSOUTN
WpWtSx4YfXQhaaRuD9azeiDxVBay7bcFW0eEuI+c/ykue02mC35ty2KOGi2iviqm
9O1947+Ifz9+R/JKS8aycRqVu1xP0GSUEIm+dss46aeNETQldTyO081evwMZ4uEx
O87KQVnhe7EXoqQ0+uug4lUE6lzzwmg/T9zPOPT7zjaxlvX2bCzJqUYUmrbejvgk
9C8QdVFTkII7qufnfMUH+fyQo18wzOXwnROURQqr6OY7Pj9A331h3gN1qRmx9RIO
PJDj+dpLjBgnqeOKZ6K/9Q092nX/M1Lzhl5vu8MPXOEEi2F+f1An9hcrMybZV9Dm
TsEt+3T3j+5aI++vlnqAmnnfdImxJJC7rHeCI3ryqKHM1/WQmpDjr25FoP8374uz
qTGZSNZx5fe16MyYSqxJPtu/pcVO1RoeIk9Z6ozk3Gk9CSxarblYDHdPXNT0akpf
kwuWImkS/GowaGLwrigR+bXxItiZIRB0M76eZX05kTfPFkqpL0P/tQzhkMw24waO
nduB9MNdAeOXjzIorX54t9u4lp2p04pn8RVgapRHEQhTge7EX7H7xPNtTtOV7Xuv
JpvPRGytJUI/p9dGdcRPIen1vQEBt+sfCM37WfaxJoWreDalocmqooww1pj1/DMa
F7aJhhd/PFjuFBRlYFfWcCWkdhErwRMwG/2p7rnSMCRmhrXzLDD7r8tA0HOiWuKE
GniJYiJZSascU5sswDnePgWeIhIW+1eVWA4tKsFhO5DwUC1AujwOCwJzTDIdxgZT
aucwo/4A6juUSqFf6vdNjb0i8rjYdGUaXl3opW2XCEsiKOjiHNDpDvZ5lU3k12RX
PowyePdvqT8NLV9lLEnVIGTCBqPaBkvlRBlF1lxvdGHdnLrAOqo9wZwCp2RZjGof
DQdprmBzUZz2efUCXtzk6rXx0gEFf1A6VgBUMuf7H+W3AA5dbU3DQW2TzDO/MEnR
lebh1LF3iAfNdhykzVc3eCAaJb+jVIgIiUhW8hIQbuI1CVNz7MPnYmNe7dhWWW9A
94RX0/ryMZuaaQqbAgpfWxZhWOcKHE+bTRBfCWn0vanVKm7LY1IG8Qs6ABzktPvQ
HsM73Cspq2FoJQID268t9CnW4YO03qBxOLZ1ei/SyhYmZvOoUdRexhuxAV7WHROB
Fk+BHUEnzC0gZy79wI+kCC7copn69Fy2MLY1dIp2m/KmAXXH5FiquOzQoxhf75dZ
cNi4+yUFpG8gW4tvfQjmvMLe7ecrhX5u4VU234pqXP3FksAQy6wWdpcEyA+jYAVj
H14X1hOGh7rnto/0Q7YGJB4nR7rnpjK3QEAvxJuJHcow2yFsNkb3hwbd/GRqCUMV
i7OjoA5FmyOk2f+aOLs+VOydd1w28NilljcTReOeGnAHgxNZ2w7BkfmBADSZu0Fi
48lYTFOw+zah7lOVEfGLAXwL9tmch7eTFSXlP7+8C3MUeVizfQrEuU1x3l+CF0w1
GXLFvWx3pSMiu/0TvYIQb9RN0U85oomU2M87ahNBcrIfz4xkLyilZtF6Q88FPonf
uU9FiHLwapLr1SP/fxw8JQP+yujme04/DAk/4wLbXCMooQWzGI7wncsHuNTrslIc
9C/oivZWnyb0wqIdbdMwg31s5iGIlpgkfQjpv4dDry32zg9vf7mx6d4rEEb2okgS
8oKiKFp2U0F8dsi2G0ANs5Bn9Y4F0/B9DRz9rvb8Apt5B6Mc1WmLpB6Cc98DAU+5
AXSIKODRerRSHpSnzj2bu++U6QSbV6bYaFGMhsPHHQl/bWXV1IRKdV1um2hmu2TD
i9svhSMwWPKnVZMNXu+tUt0K7lrPpX277JzlBUetHs5PcisNYS5PaXAb0LGV5H/t
qXjh/ou66tPl3ybKcRbjyJmbOAlQqx9+vnYxJVvFEMW++ka7gbAsLF+UCTRK8xlX
9g2XPIJE2yzdqkl8M8wnQpBGbLmZb/C4gm0+Y4mR6yUmv/bKKKM1eCpYMw16nHDD
si6vgZpTjMvBcdrbc6J2qSv5TocxDumHjfg7+GZxNso7D5AbZlshEvvwAGY7dNKz
kISp927tYD7xwwbrV1a+zDvfsDHOE6m6AciC5bmHYHs7xEWbgK4RO+Gaj5FmmU3/
v2Mt9SW7TES9NtFFWjzs4cD/gb8eyh15NgcJJnb+YjAhE/V6F1oPUl1kAPVpRzcf
O636gWMDas8Yshu2ypBCkpzxlaxtD69ZSmvnD5fQMVBBc1qJ/OY739ELGJ0wT1d0
lIyilJ0JQ5q67jA9NjZOlcBd5FIbp2G9emWIKq3kocBIV8KnZcf3y21HcfVktdvJ
B9zp/GwdOFM4PvARPagPUfYmYSf3gdIMRv0UmV4ZWAfD2iTKE7NxU8K5iQhTPuqM
Z0DLVT+fo4Psd4c8tTDzK5+flOxj7gcC/Z1P7/6kSgEiuPi4h8P9JP/kXidNwaPz
iC+NtpN8/BpF8JjIRI//BagJxPhrj5ktuoi0ngHLo46wWYjpA10+37EYgZl0KyHC
I+j6CmSLymzHhOEbhXLB7IYEoM6ehbYlGVtsBjOSJ2u1C0jw5+b8FMcsvvKKsTOZ
jM7Kz+Dc+BF0Eisdflwc/l4e7o8Nv+BMeDjZH95aIRomNAtUqLIslb3hlQlpgn/w
/UqRNRFimq91QKBLP2Ey1+oghHrZf07rUi/YQZoSkqVV7mhQcK4yT7eaBwbAp9aX
Ww0Y2KnOrBrAGJeYIqSaCCfKtgA6tblkqribFlrQ0QLEo9D3WFCO+KqMKXMX35Bh
SDxTcWYasRjolXVEQxHytMl01ojQzNdMjNiFBtZPcwOnFyWUjpGEL1A7LpuAeFyl
YXgR4n4rMlZ8/COpQKRxmYS4Nt55OxZVT5FcmGjEdFV/pvcevJR7ythu6HHXY+ZJ
KxVgq84VAxp92Mhg20yPEqy5Lx+64dj42kAFDsHlq7PLZ2GBid/ixzEIWPJyvJxU
m2iK7/EOTWfwLvCLCBHethPNKUSapTVqjfDc8qoE4wo/oMeAKU6XGmLCpdIB+3f6
u2sU/qM9KNc2zWTxVLlVePj3JbNl/aswZ3yVI2H94dT5rVhL06uJD7wmrtZM3E/1
+L1SVAt9qulyB1NtIQoDPILavwQmJrv4lt98+NkbZI3hpvWa1pTTg26kvzve2Zcx
KQmiuQS598qXjNK1pc65DLD+Dx3Se2ZsPyugLUUDhoT5Z42ZuewTjm5xJtJ2WKeB
ytloJXlA7vL1H4iuliKuN4i9eXck58Andow6B5g4qo6Bo2M/j8ovkV/tYKKN4E4r
nQQqD6zDqbiVLdvuANkK//IUqAheAh/cMn4UVjvTxVQFiho9lnyoLVLIUj1mZ9QM
IxQFKEmHa+eiQi/PtbF8On55QPGOEiHRPvv0WcAWvI0m6h/uasjIzGSzTNUviTQi
ksM32aZ/kB9qyh0FaQqeJWjAxayW/sq5vUWy0EtROFc6X4DYA+o64TzaVBbacA9Z
c7cjTwvU4Sfimy4JuRLI92B5bkyRkS7BxsWAGIsFoQKqp8DXsIVq7W8QItjBM/ev
OCBnVWsnzEik3/ZXCZgLmABsQz6g/Fp8LHfgKPjHLvRsnJVTp75VUeNv0DFcQZDJ
sVlhLDbafZGi2HmFegNC5/X9tZKhunMCid3WXcU+4DgvCZYya90xRtsg499KY4Nc
/regG/vQUEQe3T0Vt6wEQXy1Fs+K4KElHX606R3LRckAsce+wqFe8HULSjlDGz7p
OOB7VZ8FXQxKSyzdoTCHLSiubUm6A4WLPspTXICpq/htjYVReXEXQse1Azh5I9QC
d6RbAfxepZXt3A+yn6V4IyXnni3qDp4RrZfBPE8c/E/x3TE6snDr3abw0enieqXn
wD4eB4e8H6TppmPiAFSwM9nQ5GkCBypop0y/D9wifuqKXlKR9wOQJjPMbADLbWOL
Q8aekvZVTyKwuQnHHEG+nm46sQGu7OsW9/cgfDLqhjefUjke1eti0/XCnyb+uIK/
zSsDqaQJFucwveOKMtdPov8Qv7YlwUpL31rZsjQH+VzPc5N7ovUW79KLpeOiMdVj
ULvSfXSmTJ+ru3UpikY3JNM34gkMiuBUtt5SLgcB6yyQxTzfTC4EcGl8MfqfjQa5
idVqRsrTzPDBKXVCwNt6orLbjPyahW+zXkubOupUlKqFoG5f4+sSzEFSaT1e6BRI
IBQWmKlBAItmI3tEd7lkmV4Yw6KDTiTz7astaPnU0LZPHI3sJHejEhA2q+Hs6X3E
+33ITWrc3gtCcSencXdFSVG4HIyFTjJ/QWuPQ0DHhchAJNfYTZ184LyR/hBlp1Y9
xo9qFkbQVLVFYTRIhPtzfKLm7U5AqA7sMqfAqKGWlcSzLkC4KeczNIR1t0rxoAOR
GRXHacnurPGfqYIGoqjvAhTmVw1pbQtaMPzdLcDrqBAAJMA0pxhW4pdJC4oCQxTy
EuDjhFqHnrxWNAM2DBC1E1xSwEwFwuMKTlRkUpy3l9NKC3p3GmSlXdf/Bxp8PJnE
/f35WTuFqAr23EEkr5SvgcNPtKO+XVo7mZje/CpTPW6TazMmqzMR9/ahGvEAEi51
zT52CasxLdheUIdb4aod5/ztMR/I4KZ3lAn6th/3JR96CbI7/C5aYUYlJSQUh8UI
RrNWg8SvMvHz+vOjtBRkvYJL/9f/jWezjgJq0SavGITc2jAoRHjvCzJDl/yuRJoZ
DuroVC5MrkGZ0pZ3M2AkOqnoEAfmgG3jrpjIDUUAWAeSFC6n6Q1Sfp51dVS6DFGK
Q5LfOx2zB8wJwPzIpuyHZZQ0B4JOxMPM73EQG2+darRYZTS+DWpJ1I/ulOXD2kbq
n45k1iXs0UQBpwFZlzFsk+2HzCNwsTgXqsgZTztDhgq8oBRr+Vd5iFSF2aRFIHMQ
QE1wnJqcY2LczMfK7UnYF5Ef1Wi+pa20XiVPIl6ArI5MDA47bQ3RP+QqHdTiOyZ6
+yIDNBFb081Sor6P5JZxFdgaF9tIhNMWyyBHcRW5mp2DI3WbgoOxgsneeR/itqCL
oMeLo0X5lt3lRTV35BxiO4kZSeRdKDWGv1E5Zq7iHn2lWWNa58J2WjTBH+3Wmt0x
r+wwP01z1PrCl6zOLr4fD5VZ1wB63xtynLBwVApYZpDQlj24AzW4eCUSFmpqxqCE
5hd5Hx13bpGuUlavcjF3PLRumeyVALus3Ox56KdBT5bpNV58nB2NQjGgTodbBwsE
b4Ms/lhifaXmAH+5XTEkDjYVUHorxzRpkZUzkV+PMBIsWz/pwaYjM5LZG4GpVuPs
e8atT+7BXwGTMecp/PZZGNpWh+kx8Wh2IOEpQYF0DNREs0fSJaR7yyNArz8jP8oU
cJax0+MGYAmAMiYFUJqKjd94GCfDVZMJaluSH1g5OanQvPo4mvZDhlJ7bVaWnkdU
v82UkRv0S2b+reHODhYS+KAW3mH3mQ9YA3b1nIpbh6Rz6vGOgs9nFnrQRFykl5jR
qcnb62S4X2acM9rYGiqCrkMh/83yVm//7Yme1GS2zs054ccsIyhJI6Nf88Rlqo50
tQB8Ak6tMsXkhWHayyJL0h1ydwM0AZqDz57uyahpcAVlvTfDTkUTNl/UD9je2Njc
66eq5eQfqVt94tSL2k16QGx6RbOw2ig99UuL8xu2g+jMvNdrf4tzDSubIApNcOFF
/yfIc4rrJ0cC/ZqhLfRX7/J9XX6G9r86ZfgF3E0QpXaE25VW58Envpda0fJiF+UB
7VZMbphCmOMLEOvQY4iqddDvk9CkiZA5v3n9b2LotYyrOiJn4E+82nj7rp8s5jzi
t5pFZrGuITolb4SnM/PGURCJIvFtczZ1y712+vQR9KD2e6mSemH+IWViaHiFFaHF
BwwVNR9+rm7+V+Pv3dz1G+2F0RjwCijowj5aEb2pzi2+6yciq9qYjCVVJZ5uFbNq
G4hHlk0xUAZeUTu1lTeB/bBXRMRwaprHmcz4BSgwy8T+pBk88iKv0OV51q91ak5G
k0tSTqvGs0HVXp/+4dNmpkuEXv3UjjZ6Q+Nqmi1VSEpk7F0kjSS30LI0raLR49SH
EjXPkkKpp0NbIoncg8486knNLVW/Lrs5pBjumMt96IgKYfH48GTbUt8ufm/rDe0Q
Rl5vYbjCePYUcl7ZdY6kR+xNfJ34agsErZLnZhrQIbQQCXNxdYknZb0Marbl4BcY
X6fOT56Hgn7m2W1VFuJGYDw90e9/uW+YebrphmZbH9Z8YbpsltE8q38DeAKCWVy5
nGhWD2YMRXTNzEa8SRDQiE7Qs2wCfQAcJe8U6Msd4LTBZsahMLPZr0iGW++2ws5P
4f5w4qSfy1mzw7Pksro0vtp1BmhkNhGTe+zIt5EfYl4QalR7SejV06ZySc/kKBB+
Ynh1M1jMKyvoX8xIhtiqUwIWAWvL2jOsaknSp34f58UZvEfky0kxPv1/dYUWsFaJ
jeSOQymCKLhlyzKBpEO0bc8uG3ehwdC5qtGGYdUvqSYh9Io1IR/X5dnzZ8hLUEQ9
ORQ0KQkyaZhSmW2yR2Vxkj/htC+n3n9rhQdjxeltvkaleAxG3sfu28bdhkNZbV1f
i+YGSLspn7iWIFdZatbwTqmxaQUWxijHyC5Tl4Z8NizM9lOdYiM6hA59v0GLcbVd
Zzeoj5fM8UNeAr9Kl+fF2dqo8JpE/yBF2cp+K2bYy5Aaliq8EKRM85PKxMDG/1r1
LDDinBDHIAk2A3iwp7E2pTEqqoUnFm/vZL3BNrnkdJhsJIy4LEE3SFQg0RYSxw08
tnnA2V/lppWx0x/6htMaol99jxsFcZOAax/UdCHgfBB1UtVvRigyve/pBv2d/vNG
+eY9mX3lBkNnp5IclEQCJl5zITmv61u57Dp0dBGgfMyQ+2aE30PJAVQDYaqOUJU5
qAPJDepi4AtThG27mMo8zKGnBtEqPZt0nUZfT7EplfSLspx80cHnTCZygDkosz0g
T5iy6OCfPN6YfRQF+Tm/z9b8vbVbjTeXx9mE123HRjxY7ieJpfRPlI7CH1UgWM3D
mpajfRdgWqZTIhZBZsBf2LjutTXr0stnFS5txhs58gu93nhWIdjlUwW0pxPr+IZ1
/FhB5QGODMDzn+OHYCQCR6csxQj9ikZYtvLlxU+AQ/Tw84LpHfMyaNu9J1HIGNNa
KwIZPZgCS5Ox2j+OaAg/EqlHNE2WR6UfNNTjO+lqAIVSNdwnARRZuDM2kg63UDX8
uyloXTd4KIJhub1QbIKjGcU6V8fl8muj7lZlmcsHaFx+N9Kml8rqFKkOnjs/Vc+R
f99RUHC15lTvsCe4n1pbs0dImumrueAeNCai0Wv3QBgTdkdsH21oUsx/Czitb/5Z
1T4bJIz+iqZ+iVYIp/EEkyd1YEaQK8oV5ryzVVbEoUoR9wjJZRMwqG2YdiQyb+DS
07kEat07Ec3iLk13ohJJjNehkI+i9ro67n9ne0X4Jh8y7HM7TTtPxZ4b8axYHjV8
BgtZf+n4xkezvFH+KxgEgFo2y2WGulLaF5SjWj5UDTx2mDmn5lRrbY6K9iLk1c6t
6wSIJp6yNuVm2OTd6PgU3vR6KM5OXoC9Ex4YxW9lSXdCkRVvliBRYHgK8GXA78Xy
5X9F0naCoBOOT7odILLoCtStMZjg6ZpbYgkQh1IDp+Ka78a8x6GUjGB8uIXRC/Wy
DRygYCmgt0Lt1X4MK+5RR8TNkEQFBopkQaidBeQ9CUsy6elf4ukc+dkt72X03NLK
oVLQyefqOA3//dc4hphcqfKLxMr/Lb6tpJxcHlrUAaEXHfuBQzo7T0h/QFUru28L
J+Mu6lo9P5T67nA1aRm1G2OTp/08n5LU8l+YQQ3Px9TBmeiUbXZiOiNpvMKD5Xh8
8MzNARLZ083OTXgeHTYNrObWHTLH6Xr4aQeiGJjuBGf+NpzJnzvHsi2e/Sn+XsOU
95ho0UpFSWk40PQJsziu8gndchyT8T0+a041ELFaU8ar39zvFSU4RVqL2coeC/RH
bM5nlcSyyo4o08lYDAp8gnjouXbUtXzmv8b37awIo8TGC1bv1udjQDqCy5gbTtGU
sDTMfx/Ehbw9Ya3LVIDdM0h3AJAeMBPSRzbbtwKL3MxiJzBzvBwlfrbum3o+d/UC
A74AOMKThRLzCGA3cfh6NXAXA0OSs56jEVqe6xszbMRfNNWGT7rxTNdnwT6Mc2CG
LNAX8YyNrL5JyizfeVpL1JOECjF82YdO0pRrX9fgRUHW6BAAILXM8IeANVP4nJAa
zEz/7CgFNIuwCrxEiZf7LQkw2LaE9u6/R4NZh3xhnTD3BlpioAxFVelq3dE5uyGQ
z2Ae3Q/vReODqMLK5dDlJuEm8d2QMpAwXKpvtY/Ro30XcMxyjSfwk/TudVn7y1RS
xbD/gSp//N0TFTb9vcvDx9yyVllnWU0gF1SJsGpqLf/sC2fEGrFCxVVcGDx1FBwu
NzgyDRZ9Igx0gTMoT+0GAaXEPj2ifQl2iTTumS9zyeHqudAuoDni5KowLpia6egd
o2q7zkqzdFjdlwG9lWgG9fcILPrMI+x/pOKWaTEw4Rk1EQegSfl5Rb0+Y04WSpbJ
FY9sTg9HNSE3E7k9rhHbvhzeGzjOAXKex5RH2XGdN51KEw7emITx0VnEuqMKA3Qo
Rbzrsdz3bHSkbp9SxvTeuvmtDWK+5yFUS5mb+UA/oHBEYFKPxL79PPRGK5Smnz1J
XYNZnWjfjAzYK57zaqwDj/5s/BQoEO+AmeJLYUK6musDx/uFpaHl9Zx+s/bFFgt+
Jkzf6bd8JnXyf71+LQRXscddjfOwv8p8/PXW53Wu2GpLR/qaMssd5zHcZWEbPqJI
OfcqNyI8CL1BtTkI5EV8A8QtDHDZYpyCHJ4f+EUUfaXI9HKI0T/9NYFMxdS2PMn8
5z2ZYCZGHiwvRxH5BKfevVdk70C/ACOOcGK++jKqs3I/yzXSLTrnxECyJkURwwOf
9mWx7f/uvS7g0EZf0TvFBOoslinG4S5CYmYB1bCZHybbSyd0LgkVCsK+T2opRj/t
qpSNhnpzFAW2qqsgUAYr9U7YEFLe5UyJPiOF7Q0Apg3Bu36MzoDICUVf17vGZfm+
u+FvzDV3xUtr/3vbQAmQOcnDWga/qz+M2rDSdLK6XvvNEOtRwZMJDWQZVWcLEA/g
iB68tfUkH8EFhsh0ypGExg0I4sbZCpdcOU9zWrEdZ3nQoNK0moM6+0v/iCJzFglZ
jFeFcrr+AWeDIozEKM4y1+DaQToUTozsoqPa8WyPXPrWIJpNF9YipwpweiKcqAro
Vj8Ox8Z9B7ykCQ+WG/znYzEqskeXRqvs9RWt2HMczwqSe7fqvXb8Q1hfS4vupZ1m
Ct7R5WLLW/lnQ6PohG7omCh3SIVG3R8JLNYjJmkrxQgFOPaDNv1KBNMQB5+wc8DB
v3T0dZ7h0Gubg3XHpa/o5AJm6V2z2doez1bxPjPHuQLQY8OTpvTgyI7NnauTnCDp
3mOXJV86a6T7N6Ty0Ppz0IL4UE/amh9lFeIcmTH/D4AhJsGA1+EqreiObZ4p4mVs
3K3nVkHTWYxgvCQCNPQvrfYV63G/bOe0uLKDlrk/ji8ulsh1m0WTMsp8d9807ghQ
h3xegHmjImhInXggNhUZfS3WmZwhvj/wPIHSHzO5yRXriTyaM4p2jDj5Vu3E0TkT
4zGxn2sXHFtgoTzx/JgriWHY2BkKxRJnulOFpE+f94Ld2riY0MbvxQCSFi5rlmSV
/s6GwtxSj2lqKWrZ72qm0gX8GJoLl7Tx+KbBUEmGqoJSRVFvgCEesjCNp62oxuMn
92RUeFHcXdCyqPeqlG7JJpgEeo/VmB8nboeWnOYBIu1U1jHf4JtQVJjuawvJdLro
074cdZv8KqhODxNIHWgfLGJthUxVVLii+TSmTybD9A5o0T+dBxCMllUFNYASBLme
W9wtO4BxgmeEtaYRKRz9EwbbPKFN9oOREBsV2IejdUrQNEAshM0quwkouycokr2/
1DtH+51eeuuWtB3XKCwLe84CgbiC+oc7uWXDmg5EXNpmjetfYfU5FXUFysi9WR2b
WtOsfLyDty/bW6RWn92GmUTl43uDTx8w4S75thyiEfU2EmCRn240xkfPQJLxxspd
jUuJuBW99EELhKxLkU1wQ0bnxpXkePxMLMvylvgzM5q4Lrd7+fmT2Iu+xoNAYY/J
BveFQX0GAFpCZiO7zDa+w4L1fIGxm/5/A2jZN0DdF/mhEN6ybui4uF9BtYowBT7S
RzOX169IUCXWDwf15cWKfDFuivr2GVTFaWWctGezbcyByD9moseXXMFtjptye1Hc
/t+qIuTplrbEW2nSSRVdsxqNcQNqDWRIKlR3BO29TsApwqonpfhuJKO1fm5ULqv6
VjV1O5+O8eZrRqAteyYRR64KGEmiL/DXZ8s9FhTpFKqh0Slx+V+kerUTfWHEtCoK
WY/7e8ABO3U72lip+fwkb2qaMGqtfNMqj2jwTQuQkHR915J/1iY/bQjeuBXl6Etb
xbW/t4veyxzAnYF4316ldDWmYEVYDCmM3CizLWGY9yMRH7FxOwTCqnX9Z8Vs3I8H
qfSibxxP0NOjLfbzFpWUNB0HkwRorzUCLYNL3m2RkmwDSV/PH6qgpZCFFey9jPbY
IbjZMUjXjmEydLNRLYZwVdXCjzEAIFdO96NJKDkwSkneKLFWFlawq1bB8MeOrqyd
laxC0LjAus4EZlY0prsWaMQSDy5usN68OfOy96uaCwBjXXXWGIbykAFsiFJ1V1K9
81mPFZtrcKCIx/x2rHHr7MiiWAzIAD7EE2kIn3jjzSm6ZuDg7kQfniQwOFBX+0MZ
lzyutCrMKIddvXXV6cxXZP2eVS/g9m9YKGRetjO1Z7bhozUQKNETFy2lEla+bQV8
PErVWsUf/dYkQStCkzteHJUrxO4JEbvbrsku92BuUcoWVgXhjVS2MAVYOlcpu265
zD9S1RasvVoZalv6Y9rgHNAZqcZvgMPOndme8hFIU0mRQ66p3GQpIts1mwFqR4WW
Y1DlYue/L1doCba+xZgl8PY/JCdEbQdkd52h/vynzZoOBdoi0NGG/2fLXMQ7bx08
liJ6+HZt7ivHSzc1fQ2Tr1HCtH0bhGtD6oeQoxmlrwIIvJ/JBtiXlViE8Y8db84q
Q6tCoUAHKsfPedslfuGJ1qntOYcKsJ4oqcV85i6rlBoHmTlQHrTx/KV5janScDlT
zC7PFp6P7zIoKY45kmfof44+x0TjhPzK8qrcA7dOcD+GN6L7yjbtvoQeaNTyB1E4
bEvUPuMDDmVAXvNumQ1EfCHQQcqeV8YvvMVcns7zty8jrEt/d0QrKWWFVOl2L1n2
6RdqE1P+agEiKxOaFkaI3mn+H70kfsh6EdEUe7Dinuv/P6beOxOGTdTETOc+nEk7
wTIcC2FgmAtU7MPscRYnxLzzV8X0KxGKBOGRwLRjUTOq9j0PrYfItKuFoD9G7qpb
22OqnhglTwmgYWuU94ZnEHsyzyPv9cqFxHqJK5MjdSjec7Z4b7wx4BGsACtpwN+I
0h1EJQaHGilWhOv/fwoR9XBva52LvRHJT0ttiNNn0WdHzXPbAIAcjjYnYJGeic+H
IPLzvC/DQUaPQ8YMC6XcuGAZbZ3TZuwfkn69ml+mMC5Xki3lSKMMpN0GXrVzekOi
+WYN0XHKbheTeC3Dtc8fVbnfosN6kkaXiZiwBvdm62Ydqtjcu2jzELFubnjoF/ti
vLKLQiSGdZC5LgPZPQc52BbQOajamMs5RRbdAmfeC9i9pvfkpkgpCncFNmDGQH/u
LAFJkM1GBpPdu+sGvVgMHdF/WUGLWKPKR/u3SZz3C+avQfGn3fEfULNMcCbFRVIS
RV4dEJ3O2+bkYsdKm2b4ZNWaleLyD30+PMjGgTqi2ZRxtjXwAlG1zFHHodRYW21T
LzobgSQ6wFzoQmZUpLeUW6sWEetZ0B7kw5iFG6OHmWnPcr7P21p8YSzOUUPJHZpr
BCNAbaup89Mjkw07T8x/GNnGNZ76COMav8cajxTTRGmsyE0kIadrggQxwiBSNpG3
5K5+k6TQzmMCSDduXO2YCvJKZVjqM+bz0UpTksbc1Mk+RzgYLDIV/5X4uEnnroWZ
jdMuFKb8aEZPW6zHdp2GujOT1LvA5m6fHRgC78gxvZ4jimJhGOIa0VaJ/zYiWccj
NadhS259QARg4BxbVLHk+bGn74zR9BgLNV3ebxmJ+3UTpM4QoGkEeSp9HP1u4Het
LRmthqavBSknTbscuwH8QcFIDclr4w0DzRM5O0YZ1VjnTIWboWNYC+NeRAlqzqFZ
qhlScEYFLbkvRBshifj9KKtoqyaYGhHEuS4IYsyh7MGH0kWn/LfOkeka42cPRKuM
pxVfX75tG+nHW4k9y4MXSGpoqL18aHYU1x1u/rBSJeXvKKTfndgB+gPd4esRNs9w
zgl25DvS/AxCA/Zl/czEM2XQ2GFFApliGi/BMr2xpYLu7YlyyS1BVxsd0Xl5ht7n
jlrWQs57Krsgz7dpmfTmJ10f4HTr9VLVmMzj1F+4PYNZ+vX+BwH8pGPsdGIz+ZAY
GKBY8odl0OrUHXeEe6JFh1Bxi6Zsbad5RH5cbiF3jYPQQAIbw19NOXgXUhUsJStl
0jiEWXJ8+q3cy/9+EHCn0YKoH1ZzLkdkVlO2kj7PpQ/Wackdfpu/88HppxEHzRoG
eB91V94bdzbjAALfnB1ScupqHmC2u7jw+tWb7b4XLRBmT1gI1LU5UJmueG26G+2X
zfaAZaD8Aj2PgGNpjTh5ZNC4+H36af48Hba7HNdjoPx35l2Ks07GE4E0gjbULYzy
l0SCbxUgF9443PPeE7WXjLt+sL4YCYy8T+h/B8F6ie9qEor+jTZWgpsikbGoZVaq
tHn8KqlFBOjuXzNADvBwFcVgx3knEzBwYBSGpXbScIstxxEKzWhjrCMHk1JMna6E
6LZ5CQHTo+J3s+i0HN0Ow5xU4Cfqa42hOdJo7OgOZkYFncUuMC+EYjUWvMMo06Eu
5C/KPmvAKt6BUL5pj1lLQdjeDCuBVz11Rm69O/5wOKgt0hGWXk9+PeV5z7IJzJOO
tHTqzm4jHWYvdcz3EOPbm7EPQ9801TMIWCj+IxK3/f7+F9+NvR5INcOzmENdO7XZ
3Wi2OrM2L3mcMF7IW5cEUmZBXhBjsZGfmk5fkjvIIt/FCc7agMBZFgd99+OABzuG
6Q/yAiO48dfEhM50951NBfA0pZ1ntT7rU9wiRycGL2/i3sWolNcvlyduAkm2SaG/
/T8Z5pfSAYGH0KSX/MSuW2e0jOdP/1MplBM2sJcVAx2oECqpqbGL1/Zi0BEQW1X8
6G1B0ExV1vfT7Iea0imfOY1dWlcFc3Nv8TgudFfMjliyGuy1W9w1oxhzZAgSscW2
Jq0CKc56q1mIRGfSv0Nb+UspxGZED7TePXgg4nacOHAoghZh5kPduOXsLuSCo5sl
viiWOi4wNDY9N92JKVkaFmhJgn55PI9BYakSgCGeg0j8cSENYy8Z880rR8CG4Pef
8EuGoilCM4OpH4eTO6hteop934sUHh6qC3UVQldCuzydbN1nXF1PzJgWwQXhJa7O
/Jrm/Y6F5kg6cHXEmYkdPNBul4PktXr1epfiLrNQTzNgjQIWZvHK+uKjpA25ii0Z
IgRnOR05QB4FmLe9/m2reT4rWQ6deQMyNLwirka/DNC5kw91VLxBlHWO3g6/jBvc
gbE9+ZoZ2iTvUpAYRt0ULveYqOlc9YClSVqRdBDpJZVigIjdQR2liQbxNnDI/oAI
MTcJxxKO0Ch8A05Z7v5RDszJUJWg59ET+yJ/WsZRD+cwR0Tco+GbkMb+pECuFvUM
MPmmRuWIgA45LrGq1QsgIdblLAlPW07cKitgmre1K1zfAugCXHwKVYD8LGSUQprw
5P9B9yKpG8HG1e5G34e0WdtM/cSMiGRfaGt+8ff5VNXUXBp4SR9aIcvuZXlZNtL4
n3q+xBPJ+BRwuZF1G5jc5yP/5TmdjQWm/G136aWq8go2E7OJFiOG36TBXgw1sD0T
O8apabQD9UdcAY5jwz7oRTS5K1KFKWlaBdEjA0dSE91IuU+/GnjkDPmUVgR5mzvG
TuQ99773TFmWj7PKn//GGNTmU2dAvHwmfVohJyuU+ED9qfe7Ee2cOIJ4qhntVXIo
z0pVZnaff93Tlz47i3wVThRN8T9i3ZsfdfT9NJjV0+5CK+Ypt3ClEpmT/aHaDz3W
+iiiDXDmhY9VR07Lm+odxgGtn4PWHxzHWsIGXebPEtsUzciFY5A1Xe9DIzrLP9+g
8AzUKEkvrszrQsVmkpsbUw//6HRMDRc581HWYO5t8tMoZq8Q7lR9gWlmUSTobUEd
yXjfmJdhTB0C6XSpEaSF8UsMiN9/Nm2RVndNlLer9HZ3pKxTo49qDcjSntbUDh0Z
QfS5QGykPRsaobtNc4YrK2yeU5mrN2HJLVl70rwWBbRXn8GM70a+AScP3dDGpiQT
EM3ipLoae5tXFjjQFef8doWumKoditStsdU0aW/fheMjvB45WQJ52bL2QJXJBNGv
9hXjDBHxX0UQNm3Blk8LsCeQC2f4zJzFzCtJMpGkmYpW3x8qgsl2EOaCQQ/phOss
/acZo+PCn+S/tLWKq/ARrvaGLDqY1cnuHGAjjPAxDtWdBKtkzcavrSBf1epafMVc
+tzABqnmjPeSWH6vQ+SYWnfkWNEnGIyt/1ZvEfImY5DHYsgfFag4oSKQiTDaGSr/
98Vv7BNPtNbVaXulR+3jwA2d/Bn+SsFGOkdzqan4TInpBd8yfQc+lQKu6TLZehPf
vQUoNV2R0+3skzGeHxa/f/BtQ3yszrV5nC5rSXCQnz3IjfTYwkpkS5L+KcpoD2gy
IUjuW+oPpKgVmlB18YujOZt96RAs+4njLGSSlIP8cMPrOSf5NhcygtbZuTB9ylkJ
D/jnQkSVCBfygXYcU/+m8G3UmjjoRR+bLRLOOQv1Ibo0YgQpY9Vg7eoRG2WRmyX+
DUrsvnfId/v2Q/4XPo+SLyQv7D6skcIs/Zl5nXRg7XHw5n2OnZrnQXyGGxImjk1o
WPM9Je6YrVWetG+Rbj6TIKMBY1heDfRdl1b9DFGvRuwbjHtVmGFK9rTg4HHE2lio
PMefz9pPQSDzfFtCOn/oXB7QRYT2hrYi9Gys5Un+fMaweTwBuzWPi0nOPnROU5rX
t1GMPZ4sWRjoQ85yxSTcFYZTJZkBmUFNePLz3ZAJj5upt8ldG305nRr7BsfqO3Pj
LCp/AKerqkRX2+4mC771+IVZ2ACugwfPcFlq/9A92E+9dvL7VGK1WuUSt/1v60WD
il1DMRHSQv6yCIGcCxUbyFIR3tLzE3klDc67y7zLbe+w7cDRpMpiHv4GowfSwuHa
pAZ9glyDA8qydoRpbHASWS1rzkTbQNG4ioPSChC55mVOEGMA0pI9RhHadL8+jIRO
aVE03oEzd/Q7wghdlUK1qmm/V89BGUs2fP179xaiCIpmMRJN/8aB/YekV01cZrCI
6twsyOjcjq36jlEu3PW+jGz+s3iqMtMvENomJR0fIYS/IlcOb2lcRTUTqtfqwZv6
qXY8vVFzc8DMANk2Sgaa/k3Dsy9KAoWYk15355nDjIxvxnrNJGPgA+8qgbE5gB8/
8+Ag3kp1rnrBmikMhJRqmTKXzWTBrqny8oN3DNpouY+n6eybztPMHKNzCracq7eS
ftWFzYOX7RUbbMhrtAsj6HcGldoIl9mBY/vXPvsrOiFYSJn2bZxwQyIokFhbT/sC
u5AwiyW3saXMYY933z9qO9SZDPy7QpcTJeuNN8H9uLtkNyiBLo/vRk8RKSPv3VqW
/Q2cl8oNYYAJLaHA1eTJApy93vDnI2NR4cEfit0ypgqXfRC99VoTIHjyY7OReaA1
P1L8LUh5qU4C9hE/lIqECX5gZMLizLRigR3dGmZ6wZKyliMCTsaKFYuHxkIBkGRG
yb3ybZNyCa8nXSZxcTPYB/SgK6BZ0h/ykDhd/KkwF2vmcDOb0jFtH0MwhLPi8A3P
Ht9U6zGF8e6PQVubUkl/UzltwHYYai5F+gG2Cq2e/fgVnpygFV0D8fldhBY4wNYx
g8M1XG2UZSOgQBcmkv+e61xoiWi7SIuRgv2HJd+aIH8l4Yt/vjE60mW+gN3t0rRG
cmZWYQTefOUxMCjelSVcWiiMVEiAYybeDZddM7kYHnTrZd6hFLLh8nwOWI7BjJWM
q7D4XBm9amv6DZPbPUBTfIaKFbZa9LnKb9Dg6nHmbNy6MchjMqEOoSF26N+NUKLG
PYq7IZDm8BO0eof9IBNOoRFlIMdgDhkwiXDcFt6oLoC4Rr8Ekj81SnF8B06R3JU9
J1ZuIO6HAzTaX6W1Mnar/XsLQW+i3WUFgtdtv5lkJqv3e0w2GicuJ0hRfAhwe6if
GY2oQSIlT9ziQ7wLFndkNu9GkhRFHokOaYToOViRen76nCBE2ZDHuvaZH8k7/bqz
HVthMV0EyeE5WSV99bCRYY3Ziz+jhg6vKkGhFcGiJYqkzJO9swyftaTQ1FOM1YiU
qXChjIhnujwNM8SziMJ3AbMCBcVs9Z//MTZlCRrf44nGUYAxcUfo4OC2/IW1dA/v
5COVx2JTwtoQt9hmdJbZBaq2LJ44sS0A1LQgKq9F4klM+FIe4IzkcZuRMInkIzaJ
2stF9mb3QR1EGTWf7REMhN0LThVfQM/Oqt7VzNObFsNV97Z69HtYvwa1o66bVWOr
12z5Kd9hDy/PCgb54Iu5nGJ/SJlvlrAg+zFRWOfL2rsHVo94O+fy2dwsQwKWy6SF
JbXIaExjvpOi2hylghhcOeeuHHSYM4FdhEPFRfHUlme+Nt9Que7eYrCeaxm+TGpa
OeGyWORFveq77CxPYb7F9oPOyOKsc8l8OXufWHqOwlY9tAHYEmI2+D/KQ03PfuSf
gHA37iWcQVcSU8ePKnJMXTPLpsN5IbmmBSo1Pxuz0Km98JHv0y2vxKDJ9HuWfmUM
FXiUrnOOifARkgBVDx+Al+Tt28ufPx1rEV9ppWni0kV4rYL0OR/F2Fu3JiIqEOlB
SkEHo2M4++iQ1D1e88QV92s01Z5KFk4P6rTvk6e7nGj764FGh0daOMFCpkQFLJgg
z6M3AVI4uF906SUamxp0Baaxj5q0QV0sTqWomuWCUgdCsy1k2vxnZw5i2Qvgy0Sc
dtVX8cdXHFOhgkeFsX6jnUKtINBWLUB77mQWDP0/cYD0LJ3KODGINEffhKl/EiFd
wqtKas7tc53sNOgzOhhL57ZShZ6vbiNDlDCJc7RVoNI3VMvzLsv+xRpvfDUqkl2i
6GRrNVN9EBd61R8NL5SDxBG0hNP7B8ODo2bgqFVR4fBJSUyqhZ9H2bAyLMo5jI10
Qk8E7wmXNa9EXA+4x67Ezz51rCIqBErK7BFeu+DUpdS+rrQ88FMcC8fjwJGW2G/0
KrC9nnCUGZeziM3REZhZVoNANvDstb+3zLVvoWnqaDTe+SOEpbTlR5iaOe4Das74
mn3rh7OyGQlvxXsPc4glDdBatzZ6gJaA9f21kVE2Rtbzg7FU5r8VqS5cxJG/hVqo
NatYdnKQJoH0HYtvgwThSbFcMSPWq2xY8gRz57W784Eg48qxeJguuBLmfQJzU8Zb
S/5QS8qxX2LEp9o97T7AjuG17dRVZE+zR20Q4jRLpSyYaUXXrmD7PVlCyJ9FBDys
Ix8W5iaeSlb000LOf+S0GrMHLoQAYJkylUgDV8gaezKH+rsZuioSm/RxPeQ4hs5N
FcI+YFZyvkKD0DmxfWzAHfckpwHY/zK55a6l//jPfspHpqeQL/DbiP++Z9SiMTQy
wONjHdfQ9OlWZCxWkw7j4a9IzGbGUTfwSQOBCgNdCChpiMReAsjIfl6mIARVeU8T
Od/S2gwD353iNpSjio6uKDQ9ngVCjl0B5achBqqaYtd/RWj7M0Oip2h380dJNm88
tD0mBNORuxNFxZoqE2EIa6gBJZuKj7exe+9jjoYBFMvzlMSvu6DD/MVH8LI8KOAP
bE5HsyYhEfDcjGyV99c5J+f5xNl32PMc4c5BZBNLxW4QpnwzRVDbXFngfSmV/4EP
mrubkBR+r5+nYx1hpPM+nZB9iNNY98G472iIfptcjtkMVhlQT/eTLv4vvWHKFJWx
QTUMUx2uQg4CCoraDyMJNpALijkU5UwPdG1l3JiCg1HCdhuJHdUrApEOGuz5jKl8
rIsXQof56E5UpbJmgmb5b+wFysie0CZgwIYwxfedEOI2rNqDpKNFea5Ty+eBSJX6
OIgroZLVrNiG9F7ne98m+qwQz0ozbUvbwY9QeR/6hnvzk0wJGEOYO7EB1ZMuBw+0
ygNlyMirGtLFiHhMc9i+hjQbcGt6bYVtAJSa2M6w561YTqff3LA5s9YZx68jZMII
lF5vGf47MStOLjW4TNv+fCFsWzsRXqVCGd2LkAxnsvfq9NghKTUcJPhOBQ1EMnqN
tJaZ+64/5BwEnTIoWi/MxWAqUrpUw4zD757hduOG7eZ0pCMKXVrfdFEE6Vaiphue
+x9IWDppzo6wBpUkJubfMftEmjF8YVhn+5zLM7txsWXDaufjzwXTxLcXVw8NDtqw
9Y6lMeAcVdlwRI/S4DpKToVMaaXISmtJiz1mJJrZ4nG69SawvszOS7BkzXwqNlqj
iBxxsFniaDmYpdD+WclbQrsqDDi+PeioIjpY2NGhZM84Zxh78OLAbCDs7v6K54bI
n950N6PpWPK9mOvDpYdgidly8BD07M+3z1q5G4OF3NfX6+ElanN6XSoFvMYeVQlt
FnV3E9orCN+P8uN8+PHmDjtTwqzVLrSnNlBXIX6PB6Fk6nMW7el9HLe44pQZNKQd
Q6J7aXFY59/rnOn783y1h82k7GkMFHWI/+v0iMSQxkEAo3lZOzfgXPiFsKGJHFun
iNMhTfdJxELtp7Wvndda5oWXeU0DY4he2sqskB9Wqka+KT5Ly9wxABPHPe2hMUHQ
sVildZTeCLlIXqFuLTPTuxmWIwltg7om3JRwgwTrZXCWkhe136zarrGZUePzidC3
jHqbCBSoveHxYWyYAwhh6HmeHJn/yj0W5mUmG8PgPSGyAvwXCay8BB80q8LKmuxK
OPCJ2Q0AePU1aD7wTFcOdb4yQDe9snL8L7lJje6prZnnBFfvseUnZIQBnUYVAddJ
E5nbYVR9LHRnocQgdm0TXPQCMgFC3Vz+ch5fVFQ7Nz4LMjCA4mHQ32PVea88eBUX
WKoE2vcBBXVcq7MmTpxBculeS6QdtAGQN0qBI5FpjngT9wHHAWuRSN2gCeGl2IZW
00tuFOmodJskhjenPu1vpQ0r/ssynh9/xchcjMYUW+bsnuRWXT/MrabCv3tqhp/O
0KwGo5BAU1ts873qWZSdQWIMyeKPQY/+FzMVHJtWqOkAnuDEp3BnUFMA0q4rMFXq
NHifNxGT/LU2xc7p3djmlcAjikHMVnOgZtf0slkLnb5Ph5s54XR1sb+7pzjbgvgk
o9cpPlIZpmkTbqKXKHe1LPZ1QaKqHJwubONAZwPDB7xDZxnGkdJkXesB3SxhoKKP
8IepjtKrfg+BcXpaWcokYLZKMdxbH/T64wWlLe6++WoXMvY7rh7wVmmrYAEufJNS
Uc0YsINdRazlxRn0paigrEWDF/NxAVnp9sJMQmq20z8Ync4lRBXvKyQc7/B/NRQg
kKfV3En3SF6x7klV10HAfZczqDCfKFQXgBzjH1o0aeZcUOcCgXubvP4mKD7E3dsO
HOwYfJt2qaRzPUTL4gauJHU9L6ooaTHFPu+MT2QVRDr9/Y9sbxq90eHTZVjStSEq
yGi3uS4H7s2qOTj+fODoaI9l7YdqJ7GO8Fbjc0pqMCtpt4BeSKfZfYGgYUvotHVc
+ZJXQEzxpDnyHf/Vjk6HJgQI0sqwpaYktHNmgco1KopRGTA3Uxq9tqJTfkXLf1MO
clf0XhWLFWEVAPV3D45JRuwMiAbIJjsSI4lNpCAC3VVx0asBUHYB16QVXqWxN4M5
O37VpMyGL2vJp8aNZcme+b7/DODO25OS+irw2uG3ybHFUMuvv+K1UAiVnNq7cDxm
9xS3QL6nS9Uouz99JnTrtvj1XlNihTvMa+i4tQbnrwiPmAxSdsVi56wFvBys9Bdl
zrI28efkoknHlHLKJ1+Csn3BKdO0DacVhsKuS1/pgiBdwOvvRP/l+i110NAuHe85
YNYkKPcjaBAPpKnnRV3MCY+ITrw32rapoLcq1NEDSA33H9WnXgtF8NBHSMBEe4vQ
2jcIgT4eMwceJeGKZmYsZ1VLUq60fl+C2A8idr3dmktV14I0F4PDPH4QZiwdoFTw
WNGCuy5n5OskYKnvQ3FyaysM1ckjG1k3Hb/Z9b5ijv0GHuXUVxmocb84Xm/Y/8Th
7PRwYwjGzdYYVEKsvK40y+npl2j6Po7G6N7y9vj56GwCejPWLOK3tvVkegdmjgHX
ChW9EseO+QxfzKJ7APBjad2r6aPd8cAOLyvLEv6nkPjpCdR5oCXTZ3+5wmn4wHR6
K8DhqXifBIQ68n25VXSBVLMcVhMzUFJ/dqX6bYygJv1gwCf00VQBLijEMG9fw+V+
0ri+qZlUr+Cv4m7vyAPjCrTHCJdN9FKshEuNfsrChTrKi0RMT6gPk5wrOdBsIFx9
FH1uaFCyt6srdihVVRMI+OJmhECtypJqgal+5TdJSESW9Bkxp8no2L08KXGESlNL
CQ+38q66MXRtjfEbOQ5IdaWfVScbr9EtDpnO70H/cnHxdVgdbdCEspx93p4KnvR9
dYSt0GFraq1ga6LHy7MIkWylageJ5c4pm+1CC4ycEd9hJIFW6JOGRi3MIzkl7Lxp
SZ3FYhgJZ2HNgkLRahGM8CPX5QVywjWDP8xCWswb3athtP/ezEU8ffI8G0nzPLbV
jv0qXGS3b5V3Qf7EZl1W87hg4yh8Sw2wbxRrKX6koJXomZhQFzqE6F6119DUKxfQ
HMYjXicgyWUnY+Adc+i8nwjy3oiMuIb3X8F+F7ykGRP08UsRt5bOOpz6TiflE+dm
H1dcDLb3HOiVqVJvQZWMzKmM0/ATrxaTt+CNg83zqXYw16tObnVtcEzH/ID3Tjxk
qQ7D5kqtQXjGw0k4wQS4rRcHLDXXbZ7fe64CuQluz3iuJ23Is5umC6TuoroJ7JU4
qaeU8SQ4/NI9qHC/Ybgypgc8DPaPeFGeNOwrbNBFPZbK/TDY/jKrtur/twQxFBw/
VjYt2mP7iHldYrd/yLbhiNHOwoFXSTHKmAJuulGfdYcsWNARelG91ZyfxLoqI0Xv
IqXjiTeH4Ay7IsUBzan6dksEMVH9YbN/iZk31Wnm/nySQB+ucrkOsuNAStihkyH+
C29nWFTF5wjGIqM/jYx0H+TgAnACYbFz/nZ9uz+dxUeJOfQFpgGQjXdf7ZAeIrmX
u9f8v8FObQb1fhj66vCAsUndrsGcTdN8XNubeFcF3TSUFP16UzQLszXqH1qRCX3u
6UPIe2jbsbH7MpblsaydrlWmRR4GiMclfZfz3n6aB3ftVsDYvUkleCG7P9+ntwpu
pmeeSKRy6Dy2GIM3DLCYZOm3FIMTYZ8B6lfq7IzGFjdlfJhIdhpZXVBi2bezWOTg
X3UKpKAW0ReE4AOOO6xXVjFLKKiLv9AKnS9Yd+7YTuTo6xv8ZnlFiMWDcI1C/zhU
HTfhvsFBcotcz0gs6JlSigQNBLkceE9ff8WVt3DLgAWdDcb/maefxcraEfrS6LHs
xh2E5DgqKTMT4OV2s0lzZg5IyNL0dcVdN2712HChMUX5Yw5H6QuyRUivquWm6I0N
WkEBaNa4/nGZyVkwFAsQC6Qv3xiuPxkoajy4lAAe2zZyfUUzOH3T5F1Rx28cm84u
cKCswjsxM5elBFWL6UJcjGgCRVN+kvqHwICnhoVdtHeJr/bszkjhbXsUrV6nf1Wg
SWggUyGU08LHYoWNAXHYBNvybHMyNWzn+hoes/vbTZJCNqcC/ecRgwFqoQ0JWp59
drQqpI26sd4c0DPR46eUbmX6oBZQCyxmwPawf+wRi8QWCTg924qzjKnt9d2A9euI
xte3hjWivBm72fR8NvH0bygd8kY59cCS05rDjUskPq0fv2GhAxijmWNSzfFrY7YD
3zOoiUJZRrTEqGS3o7X0sQJztB+qySuPszU7rqEPskI54geWn9c67aSGPOoJOz5O
7spkonkCVrc40134bHlyUGYfcAjLOGJ8PsQvlbmxQ66H/t1L2X4p5ibfO+saBBbZ
fyFYhbM2F4NfgWxsaF0lQpzNWo735DOfIt8Kwmq26xNhm9/hCEXb2VibTpGvig3/
07t+wFpiuQgpwmj9rK/zfPT2OQcrHh5bZpcwXezq2gKEVX9aJr66NrqGqCSCj7V4
FpBtE9+2uyWi2hNWVWaXpZ7vSJv5N4DMAG1crLeTRSCevLTYpqoOuiEGJB/teFTK
bIMN3EhMHtGNoJa0BeWGan3xMMQK5Dn7ScxMOFjh5XXo1PJZ9fl94nqVq1FMFSeH
gwSAL2PT6cRhFLh9jpF1ciYVGk9E7H8U1OXg+ESCQZzVOCRjhsZcAupujhhjvrpZ
BiXGNTKBc6abxh9P3wEnSNomDrbE8LqxVQkS1gBgJA/NxpqIotEI8DC+tWauSdK3
cq97ZkDopZc61+ErWh2Dhyxz/O6/xEtbSbdlscKasNhD3X53RO9XuAfwjTiFekvC
VPRDp5c5OsFWYoMpa+2CUaGlVm56KaruaFyBuxaP7WlrOGoO4EbXTZHLY2rvIH9n
Vzb7iO0rzoYosNlrJ2e7O7ZDsZ5s/r9UDoz9QWlgaWteiCSyjnOipOqT78s24bKY
cpVW0scf4ayxs6p1fmvQ7/IXDugSwSYO2RHMr8IZJADzR3P+p90RFiLRcHFfFfu+
d6hc2KGY7tClJy0D0CO9+M8cFQvLEReZfI76Ordrzahzfh9ZDixDP034667DKwuL
YWMnxZPnRTg9lr2Ra/8QnBZLmaqX1QQISAzsR0a1z8UkUnKkHA9nXiGJ3BfNoMdM
hR3hkztL9UoMvN/M04rlUSb+VCFCKjo7SshyNrME9ThhV8bGt+l3ibP6wHrVVhQw
19Qt1xKXIswQWC+VhzKZqTLj6s3vWxZHgwlGgNpNZV3yBJ5MkxZGOSnSjRpL9ygX
48f7KSZqhNd7Wt7ex4aDXFnH+lyjgxkNsZ+jFkVGRK8opCfHFEzyjfH6WYd8d1Um
PSJs7dpimsV7PmutShkdiqpvZDxi+oxA2cyd4aH6jF1wOhSVP5OKpyEx0z48K7jz
dUKZg6xrk6xmb/UevyALaHlOJyVf7u3ETPekCA1wUErrytZV4fRrpbxeaOL1p2a+
7zQDHNhb6ETfzbsniwv6fhM3NjGRdx39kFCukVVCMXZKqaGvVTQpnMPo+DftsnlY
5b54b1NGk6vut5CJ8vYumjltn+MnaXt+NT7Y9HARjZGtz6mF4QVNayZRdpiXZNLk
GtKwDDRLDJABtOHmacr/LqcJT9b6tOYEnaDSY6cdnlnk1DDQm9rurtJtP1IfFSM9
UORTlidDIKbqW3ygQVSMW27yxj03neCi7vOH7hvA4wX1NEiokj/Stkk8q4/JlMyU
GbhCB1qyGm1qv3lblSmRlqASZ4enC61fHDMY6k7M/35QOfWhlmwhvt46U7SL0pvN
l6MoHF4j6Yc8Tm3u2UxjpnfdNiECihNSWMx1WIT0JsoKYkOb6IcUjnhdtzIRji+Y
HaLUlzI0bRoloN4DI3etPTjHoPWQ+lpwC55KzKQpF8fcm1lJiiJpeAzz7UKqIWxc
Su3xhZUjU54tqKize6t+yfL1IDsDDqZ46/9H4ZTivgWrcB2973iVnrezPdmK/g6R
WOTLvCgMXNPo3G8Aqpj8Wv6x+Kpa1lP3+n5xcoDC8I6pkFfxF+HiG4DcoDmf3NXi
mr5w21uj0bWFTxJTuOwUNvrC5PPWqBuxOJMakuOWmRoPfWepaMvUCXR542oAX1wj
oAE7wASdowgOxAu8iFOKIV5H82eBaYN0ZNd38r6caJPev2LsnmG15Z87sMInuwud
zvfpC2p6XniZW1sLYVIIMutIba2raPrAoaKbOvncDb8Gigh76hEh9REXj81SoZRf
pAz2dw7Dw+tOLvAAD4WI+VkcPC0XF8/u4v3CNxelT5I/TP1WhP6wOLoaYNpri3JG
qmuNxJGde56j2J/jfoOBGIU49/+lJcsp6N5iTDjcukkWSUzJJZJ06G2IDWz3t9qm
mYv8eLf07+w58pvcsJA6kTc7f+NnPkCm1SReuC3T3td2lV3RL/6tFcyQIJxIfjKU
hmX1kpUyzwLQQR0km+cpNSp7X/9qhwZOzJNXnF3RKbJgPq5Www255EbhAICNSBb4
J6X4TgcRYxrMIZ36fDrKZvEVWnp3SqzB1ZPVjBHRByNyR+Sl614McOOIGGaK7jkK
BKEATi1YzrYDbnZtJPWBmhPaBgqEecPGNTDPjgxgZu58dL4HkHbal9Gbs36d7WPD
xf5HOpE188oBeGqaoQSTRN5ciPHgZsi6fMSZP/GHiEcZLUEP3nA4Tomng/qzwdwD
ZwNiuZAb9z1oBrf4tL58g1aLZRbK2z2MnhQXfLKnNRFFatHQFg2ZJg4eCzx4ksvp
CFBVHDMFStRouLMCVAmg8Op6Jresa+/3xmrqkmtl+LKWDWRi+ykdz+zO9+DhybZO
gMdYhJpmFqnFAGU9ohidoV/IjjEBhrf+A1tA/y7N6mPEwbsSlxlNNH6O4Gq7RSgz
UpNJvahdoKbZw2AYE9gZ3c09NYTys7DfriILOovNvI3nrPWqq7EH9Gd6R+ze3VfR
DzpQm86MIS3FMKlpwisFMFHAwQYwUd5spYn9Ju8ph/KRiORDW3j/bOiuyu36Iewv
/S/qhN3dUTk+PIpe/v/lp6NA4CLVqd63tEitDo96Zl9rYp+fGv0fIv9/k0PXAfKT
XjudxVp8UOby5K6g+NujEVVjDytiGkHfn/gnKo8GecdZj23HC7Wk4qKe1TZMvyb4
7L/B4xFGcc/xYD/tEyy6jTR4F/buY4jBNGBLsT3CPNcUAl1q22Eat06CJDt6uSqv
WzBORWEBUO6219y8kmaKzTNaoGQ8xBRWb78rUmsMa3FTnUPrwK1GC3FT3MkzejPU
m6djIZtmFASRwrYXY+zRWhd+UOwGjz23tpkfUh4RduHQ5OtnzxYf5NLNYkxkcRgg
MNcbhCXaUlgqmO5b7yTsKQqQpSm4yuyqQo3pkM7TCSajq/oEHKmXSkOxknMrR6sR
He5x/1pwymWJx9fXMhv5nsus4kSmEcOMF3LhLdiCAh16DVc8OBPqkL5J+e2uU6qD
Gfh9cganoA5w/Gvqz+qJ/FetrmQCRuxmv4WJZ4/LEmnNkvBrH+gf4ysLKGW7jQiF
PFrJnvOdgPPgVEhSidJrHMIvk/rEuo4znlLigfdU0VHYYt34+eGX2nHanOdnU6eX
hqI4hFm5l9OmcxwMOlbQi3QtuA7NtX2hsl4vncxH4m93zDc7oDA/VHoRMgAFdTvV
B71nhi0xMfBAzR0Cx8D7ndas72LyIc7YMMav7CqhOzLAclbVYTMz7zSmk9aXcqiP
KLM4PHwxe8lEjlmggeAM2V9uqCpVXtyOlDgC0T+t6plgPQo7dtwRfTkzIsi+JfeE
sHj0G7vG7kyTwHnFXEICr4L2/+acOkvhz/1x5MMdwAmZsffs0PpmikmAqXzLDCca
JSJfBnLCtCPGl0XAabxI+ZIc1Rov7wnsYhFMj1Jb0+yleGn4wROEtEM0i8xp5UJR
VCyfspFcgJM0TzdYGW4VQbaRfWTMiwpr68XVkw6cPa4CcEsm22DxJfksbGYU4dtB
AqVlodCEA6SOaZ7sEU4kQKPSTcCbEoU3qXDCCiN1cbh8fLGqHGj5xPnIWTHMYze6
hs5Y6UH/lbsFp3ywCQucCOgkkJjNq79tvcvzNFM4z0bgscLkDVOjRQBSITlsEQUh
/NPoAW3bgVq2q468z4s6tqxWpdIaQ0fs79CAEp1QIZ05ahqPcPC8IWMP0u8mTSgx
Nx4kog0R5yOpmm107mEkgsBWqDM1JVW+I4SEzx2H9JtnPo8qdBsdSQqViYxb14hF
j7yU716CmYUB+aRgtz95px2jwZ1HVJa4JTuzCPvOu67pyLtnU9LX021+gBAfutjs
tHjQnsTwqrSdXbRmnQCKamIoMvmqaqtKxeehjMSb+vBDjU1Y0iW93/I2kvH3CBtu
TJm/ZfR21aMRSzNpcISk4BXnkdtAReFxpXPbSfpJzcgmiRFnMgj+dm6MCMzD+cbd
Op3q8MM1c/MDWG7j5kTqfx2HhQvGIJAPqxe4inx6KdLs2Ytht5R2l2IiOiltrm8w
XGIp2cPo0djHTGQ/Lv/rk01Cclr5hvJ/uyrq79kSujsfYmeq8Dsl6BF0YYGOxhVj
F9bsxHurcxCCssM3yR+58J+FAsUR2Nl0ql4EX40CiNOmDOzP5sybPjiWMfxuVjyN
2TuniaWPLEb9gDFIxELnrp1B5CP8ICizznRG0nL1xYZ2VtJrIC0wZ1lh1RXnUn0m
R2aJllTJlNGE07G4wAJtGkvx7W8PSgToXIGnxlkZ9vAKlT8HzJt5ftEr8rqkZUFW
Y7+HZWFRMAWk2JNQ/GCE6iXwE0LrTa3aIpEWCsIHsTDNx7oPKEKj312qtp49MAC6
qUAhSEF7AN+Rs7wvACJPXTT/R+6/KQ3L5lt83wjxmJ8W9nQtOEKKbSAPR6B59UK7
4/9RrKzppLPnYqmLCUZV0ZLpehD1su5nFxA9uxn1pY5AqMoitQy0MrSxjz+IHwIf
k+a6d+WjzmHocHaxoEKeXrIyIwInByExi3i9Easf9T50dy8A2UwPBSggghRe+ae1
/u0578yVzRFu+q6bzReRwPfLeABqH/DJedP3KITvQ1AT9rmghikm1kMTHw7qoOlw
7maE/xPcl2OAF2ZPiaBbWcA3n82sakVW+6NeMx6eETH0i+i9jbf4WMX1ia5sIHEa
79ODYLkS11te4weRZ6vLenHgcaARgetH1E600FlIpKt+T7o5m2T8tBA6Uu2CTM90
upt6HAITqhOKxMSnItFYVNjSM9l21R2rWQpC4qrcy7dCJsSHAP2o4rKeiUu+Dm5Y
GvAAJM7y1ClBWATr8C+RfFZW9DhEHQL9wQ2F3xZhW7dIceAfMbwCnkOEC36RTx8S
nni5w5LHF6LG1EwIWtYTKSJ1RWfi8KZFdfil1ANbjpdebX962RiE9zoPQ7iBs7rI
Spnzped8btHnl4E9WeAGnhW/GH6dcuE48UVczR3WzivRL0/DWnjqgDBEDrGBt0Hz
nDkyXIRf3q7y0NZDKQos04eGr9M9+KQIZL52LbHpEeA5QUOnMkoBfXPYoB+5fH4u
5IJFObIo9AY6CCkY4JMhNFLNSHXIr0M/lQOZI1FockI14ykXWDhm9e/mBOiGuVqD
QOylbtEXCLf/bt8mxDPHHa+XZnsZG/JToDywONKRhG8FqqddLGkG5EOwoT9GZK3o
o/DTIvEqNV71DjT7dQT+aIRsp/RT7wCJyEqRKfws1f4IkCIdKQkGkDasW55xD0v9
hqukz93YFr+2h2go46RvnfhGqE/mdrkI3DXMb00W5BbVeRgK7h2liIzKzmpWrcZ0
54Vl+2WUKgdb2VUozBT3MdpC6TFBBT1XMYYaXonMLv8Ev7kfLw7Yiqwwcv06Q6KN
R4NFowo8jExPwzNa/GAUQUlqtHvQrnx4wW51pHmr0pRC+7wkkse1B+2GAyIlJDaJ
wIz1fSHcNnujWpFHVAG635OLbfF8kird2wQZOb7Nrt8aIAKccRtLCd6xoaVqCG4u
EKkyp6riKmgOizakV6EaYnxJTS7KE+FjQCrLBntve9pHmVvzAqD7XGy1jUR2sKhJ
pUtx1IXHr42Zf2SfnVXNmM1Eq+D1XJWyQ0EiaWRJaKl6HfvsWomgjaEGhdb18lwS
vWEATy6rkLHQhruQOBp/7K9xZ6BBpaDRKfhf0WAfqZsKHMDHVc5NTPaGNd+QICd8
1068A52dbC0eDdVxSgrpJVCoudwqLuMweZkDFAeId7cjxFKBtEiUpitYuaQI6iRG
4O8QYspFtV/OHouYTrOyLd46P+SL3Uoy8e9VAKTbBx5OJZ64ABusyNqII0Uz5iz+
h/epcFufmRitFCzhikYHPnzs4t/8s3+P4O4EOopuEII943RdUhRYfLglojzgU6Ac
YNvDYsZQwK+oYoW0yA4GYkXVXQJtLngBVD0Kd3synGDeheKZzFZ9Ls8IMnavW79J
Q/ZAR8wjKzRHk3voSq1Tg4jixl+8kFyii2jTdyYQL6daWJIb/aUuAxeG/7RDmmVM
ElzzD+fPd+MNoCuaQ8m2QDfLzQAXOf6BdWBYkWMkpAhXU5iQO5WldwH+j1myFlZ8
JePuXrvcMSRb+/5ebgh82gEn7cJ/so8e7mwc1G/U4Si6KD+XZd6kegGNc41mFLwU
htrtdqIBjCZ6nVh4NqY+d2nc6llzuh+EcExs2vRwqGBlcLOMCMGYe3rBy6sAX9Hn
CFp222qfVMvzyHS++lmXJMB+awY2eXiaQ/9xg6/rtZfzlIgaJpu+l1kqQdqfBEth
fdvJP7kht8MZLskniJ/Zjhf4hckPC3+q+JnSaikrq7pSR6tKq/KJWDUkl6jtz3yc
YCkoEKCE3/WUzDfVsWI+apkYVyqHvo2Bi+4VGuAyywQsOIgttpRWXEjzwr4uVGg+
0P5mRJG3+/8QuqQrv7T9JMrLgVhP6RFwhO01YAhWAuOd9cnZYuyAuYo0IXCtfqca
s0kdO3MNVVNM/YrUnX49N5SWuZlZBgsME74PkAmORpByNSsaJDKNoJYe1tKzv3QD
oXnTRILxlesPR4HDX0Xa96odpKOOSRDbcHSjbhE/RQdDT1vUy6xDcN23qLE7R3XV
OvExcvnag3YDMrYYxFUCvmNaXrD4flSsKkT7sei1vOfbRgev9NZADDwojVn/EZK2
8aImEDHf99DWmh+K2YAebPwBKW0fkVrk/YPumVAiahBDhCa3djLYQ+O9E6LGXDKZ
3An2smiwBVQ48MXtr9w6INQ6yJ0Z4lPn1kIIQfcZaKivK2WRoMoeukk9KOhW4aN+
EVW7i7+a7Sl+EJQFVgCcjArGfNWYnqnEaLCs2QQ0u6E72NlqxPeUZFbKLsLexXxd
avLeLrBgo+HN32XuLg2uUa1Xf8mVa0+pwLeoX1BZiRdXocy0AccIqNdCExmkoVxI
wp4wFb9RV3bXPiOhx7ICDa1XBVAdbsvifyzGkYtIxw070ocI7HSABrYyWxgka2sv
sQkdjJ+KW/Isx2+8jtVV4k1Zqlj2VXo6lREBfZ/4dF8Kx6IlQ1dBSVAVQpgg2OHL
lhFA7Zjlov3G3j7ZPBDot5nGe2w/qAN4sqqBC84NmJpWp43yM4VSNHLGdHDXu2Tv
Gaj4llE5mQCHB7GEXuCaEzwWuAu93VqAJcqTzheLTiGlRK7X5I6sbDp5Ua93jthy
Uhrw9BuRTR1nhW31uDDJMPzQtoEorzlLX7GCOctrgTqQmyfXXtI8EK8GvT7+zIJi
ot8bGINMfgo3yRhEYhR0kmSAOTVIk4WmBzyvLhA88a8jVrph2Cw+v5p2jNFZRMi2
XGXX4IfGN4Gk5/QCgdPkbRoe0r5Wj66Vq9d8h5WwwYeQJ+63pxFbmBBEHDvTsMZ2
xPBaCXZSanY07UPcK4PpUP6V0vCaU8gunjPFxbz3XAr6bWkHoYMC+43JjSQECjrc
rcDEW8Rqc6Rma1f9vH0BYicpnRTt0fTuy9fWYpBYsBBD9d73E5SLPex0ItTE4k5m
nlDRtDyEk10d3DeJQhla9ITKthFQocj8LNycac6Iv2xTG6tX4/ifidYXdx20uNkk
sLCBqS03OkS2en1VOGM2iTS3hkI24LllfRRPQaIrFR0ei4Mg0IaNJipCEdacowfx
LbdVw6dUCSjfw/zRKXoncBOnMRZfyMhH02BBiV3wQzqEETyhqXsJhe/uMNO0WQHb
/A8qnAQba0YnGaHCcNqvgPR0j4HDX06fXZnIXBZJRM8F8Tn9HjFhdFiyVgNexnPP
cq7IH6ICWM/1gNCLfVfZQCUUnkAvLjjxnoDxEFZjHk/1LFb6zrfwBG7LcJtdJ6n/
HJXdX/6j4L6ePfOrA360ACPZYDnSp0glh6kZS5H+gHERQCj8OIQwAGrDV8kn22Ao
00MituCo8nMzk3eKeJs6mTGqGeWlJVbeYk2WQsxhJy4zfy4kRMTAdHKIYd2Vq3X+
gPzPWrst79yq0ZixvHBwAnBYuFk0uyn5Xd5ST4rQoTKwhgphXQ4rrsNO/qBvMD+x
RdtDJ32nUJ/aocfwFNKXHna7sP4XilIafp4qMYqHcNGhAVr6dSi5PxiS9tIR5vXz
LqSmgJWYdMMNZS1qj0Igq5q454tNsD9lmFxUPLb//EbX92cWRl+uSI86ebC8fc6S
37WXVIaiypiiRwrYZD35Owt2xO5t3sXgV3wONp2429xpYxZG0dIK5RFKN1Ya1ChA
tQRRz36PF0hCm+b5+eMMZ207q7cRie0hcMqXAjyetarD5sHh6V0ucHaLzn6v7NHq
0z01oiD1cSxhwgjEBzUZNoSOdaUlxiR44U8e1fOoTE40q+a4v7G5rA4n/q9HiAgz
8r0CttpIRRkRr3AKCUsaOwLSqaQIql6yfsWg3JOtpt0URfYvBG6HKSaMYz+6+q6g
1O+tVFfWJd+74vYLuBv976oy68FK620USYvGCGU8V020zvLaG9gXT7wo7FCcxrVW
i0TdEdAvsOKM3GXQywR7wXnO7RpT/9r9+R/SRG6U8QjmB6KXMqpOd+SFwbCDClUg
g/dr1J6AH98qzxgsH5MtytiImS2Wd9H/drL19wWTejL6OKkOkOHK8CoFz1Px+k/A
RfNkf/ymnn3NKJBka06pe3fwiY5ztVE7Ptfv0s9WiNm/cQ/rsdGtVOJgrw+1yzrE
B/1tIuty1z+ZoPBZSty0LIYm1Z2x5SjnneuaxR95JczHCclwprl3Re1K6+YRzwRU
ArOsHmoPwt6kg+CN3NVO+q9Cjpc8dJ5ow/sNMWmSF1m4SWH4bDFUF/r3j3Edtjgb
wHiONbR4HZxHFEhAZuCH2UvZaZLxvlMGS8CBzuzsrny83XqpMsktkWvyTyHaHEpY
NZPnD6U7P+UFmCbSCSZU8B1UPCco09QLasiOoruBq/JHYgxF0bHR0rTX7L0L5Hq7
Xq8J7EHakm/6jcda9hPes7aAlJXvBK7nnMDkHODee5lNfNlKhCLtUK9TKNQ052lp
Q/Q2qM3HXZj3/I/ofuDbqSFeBnSRJ/lw9WLq7GtTYYqfgmKLnsV0vdVyFJOToAE4
Docj/IITJNEiEI0959yYsZFvoZj/spq2n1nUsuaGu8wzwr/78fg/tDVb2pbKEf7w
IoLGplR6E2wXY2tBs7wfwHFDfEJ+JThzo1oyJeHX1CC09F8lRTeAOAjcPMGGLLbv
68n/DMhQ8m6AwSBh3YaQNjOEeMMfTZqocNWvVs1s0r1TD6+YNZtqnBdxjsKSEGUy
a+FS/xhVRsxfoMj1R2LsPCIN3CblkIIp4Qn+eHI0vxupACttHTIXyhWyC/FbNVn+
sr6p2j2SBUWior60FHhG/P7abRxjhwUnVbQhOzBNg55AldKMMnBQ1C+yOm65eejc
HnP/FaaLGbO636ipSlN8juu+ODf/RNK4bGRQvTnNb1o0W1ftQrCkiVlPflVSZE3U
XJ1yWRMUgvtGfozYyWS5Q28PROBpo3PLBwdie7CNR7KsdK61eI/3B2bXBc9qJn3j
Eg72tuqMHhy70bUozHDqi30LkD+naE1t9/QD7RsnOhb0OMM4c8eGIIdVBqWv3xNn
z52eMDiAdfRy4aetRfBk/H5KA1n6V5pFos2gQYPGQy4ARmFaGpPhGGoh9FCQGOdu
Vn71kjyKK9Wn70N3yqrT/F4c/5MckBgOTleVgrLoDWQgeTLn1GkwPJMB96nGdfpk
gGnmwrKkDe1gYZkZR1kp4Re7xFtgQMMPd9Aw4YxDwCMxk5THXg8RG+Q6qzW9eQ43
tBcEydylzcvSywDcEQvy0AFn391H680kWkMeHjIMrtWqPwqPzc61lIjM8RhZ0aZ3
MyTzWa1U5AQQZYQUbQ/+7sT4sSOn6Xn2gkkINfgLE3NxzM+vEB+Na0GyDoMhfoH+
gDptYy3Q9lxrTpXX2l7IzhNelyYCv+WZ4zYAMNqkAv25zcBQ3D/yE2n0W3U6KXA5
2hRqUQqyKXDr9KFIvHkb80ITHjKZC0NyhH94GtQcLgL/sgmPxORqmeUPn/jhMVxp
x7FjuzsDA4FfZXuG6OzSNxUEN4aPNZioq9bTAOw5e+k7J+Dsc2SCHl4z/LRGNJAL
0e+9dhHKlWcJwgfyk6KRYf0DDs6cncKR3mbQ7tvfoybaNnnfo4AzFGklWGsg2xvU
baL164bhqdHNTiDV3ojuBGQ9siGRsY+RdkQ/bIa1oaiVaBCds0djvulNJ/Lm0yMG
FawbhkrH1zTQBR3euCUqguDu6QGwW2rIZOIdaAjJ/gBm+EtBZy9FXq/Q7OfgWHGj
b9o3Nnbgc/6akVHAcAgaTd0VeYxf1oj2lin/caYxGNGlAAT2JXD8ddZ+JUTEI3fL
upwaXRVNLQr9631BrXzXp9EKD919J2MUnn6J+lzA9ex19nSHj6lz/uZ7LMfQjCNT
yk9OQ2h37rDzyjxPeK7YvDQ339EMNexW0She21D6++IIJAU9yab3PgaqCDOBJL1U
PgYvF1t4VvSFTDR32YU2R0iWLd5bYXCKNbqmryjOk4m2e3Isw6SZp0epKpHB5eb5
1ZLoncoszsq4rQRTDHvyWTZV/wLvMhvgPXQ9XWCH3GvJfk8GhRfh6QE7Lggqi86s
jXjAnOS9ebY8eH1F5sTckFFoJBXVtCPPkLf3j+9YBLLqlDRHUK8YMUaFmlMlpgbO
nx9kdCT0b+dk+/OI26sMrKlD8drRPDirRkks20/wFPAXz8h0XK64cmc01IAnFlUs
mt56FSYYApH9Hqz1eaDTjR4rXgHERiUuMFAUhaqZr41l4MbC81VbsiD1r2C0/TJJ
OjIn7/tAuYrvtNyyUQ7LJr0/D7Y1SFXVhYihZ5QDhej2udRV5WNhkll76Y/TEGhY
ve1CwOUeQWo6Lvl5x/vTi8UDLwOAf3Y/1AP8V9L2lcjRAS4jmxGFAytAuY3YOjkn
qqEgpayJVPE8pLoYIhfFxqvzyTUXuxpHBizbjJJOqres7uiqQESxEM4e6rSl99dJ
KlovZOzP7ktlZA2/DHh287yosXTN+zqO+4EanuMWuoyTFjHfbEPbYL4QhuQltPUm
3VWSyPYdylz+QkpxH+Vf2Q4tI7bnfkdVjDUt8pBmYB5lWGxnhzRJ+yp199mAR+CP
XxUTyFg8qbj53fisbz+ecLCAQD4Nsidy+ZZtuC1/sbGxkVIeRLE9QZOmGoLjlom6
5VhEvUzwjUvNYArxEpT1kODx2GZtbfgsOs4ANzT2J8Fx0mYZMzImO+nvRTg+iwPe
gjMQkZLO11qGcwR/3LowcBKOo2JwZRZcllwBex8ujCzmsFbCcezH+uWQfH2WJ/i5
90bJh6kpLnwc5cPMLgjEQMu/PFJNHb4814I8m5xmgI/l7EAlPEl2fcxa2r4Af+g+
2Nv2Y5QBOXbw0YCEdSrif+kjNONNSAFKOELneK1Gc9l7j5emhO6AOu5inIRyt8Tn
C60MACqkn3MRCNn2HITblXdlAFCA72QGr0S1KOS6iQUHzlp62X6T6fKtOCStGsI1
aOdDQhIRgUe457VSGuFf3lwC9XDxWaw5NJyeSsgO/+njjNDzf4+CilaoWGZDgtP9
AkDFh9HOVseXR0qLIiVLyJ1LcGH2cuSiNcGLzTtba7Wkl938kYXml1lsQyYkDicL
EWtk4jdj2J70sYznj6UGX/LIWupb3UA4rKNljLSSxMtNiudnMe895p8t7xOl1OS+
ndvdvTw5K+dj0ShLBXLdYyuQZh6T6gwtKOU0+R8AA7YQmUKHrej9XTNgL29xZWU9
UJWVuAS0xc7o6iW9kdLo7TH+Z+2RTqugHs21hoWz+WqTy9OZUkeLIdujXewi9zKI
L8eRVn5NxZErYMQqQmZGJru+rB1EHgTnk8GV6x1vbzCo/RIGkXnspJnIKxM/MtUa
0c3Vr4/Gix8aL+XhpVlzwgKLmJY/YYaqvvpvstPrbAWny7Ljp024piBB2rHbymNr
wa56WFIwyDiTC+i230mD8oPyOI0JCdXSIOHCx0SxJOvXSuSt60ETdPW+Ue3MoTs7
qibgz1Z1M9rVzllaqHadyl46eVyCnvKXyIlxV0Tm9KJcCapXd1ioOKj8IdlCWMrm
1Kr4ii7VX4ngBRLkTr5WynCDBpd2cIyGAd4Kt4BYQhL6UEGCP9lbumNWTf4gHQjU
3Gr4QhNGir+lyshP+j09aBDhJz6PIttu6HeDoyaJYs5d6REEA/CNgoEyfeKJMwlL
FCwzrj+LraUp6Q+t0UNjcoH6dXMmLtnYYR1HlrFylojQR35rMUFe7ndvjVDRFvjm
qcnvVmOXuLNzgBHUX7IhsFaTxEw1kcf5M4i7NGEfIUrPPGBVPwfhdilW1sZm5rSH
yLpue+vbDhJkvASDSpIdzOcTrAAv+Ou33w34Mr5KYMJno/Rb2/03F+u/7JoaVQes
cvT+be3OeMe48c2lnW9uFLVU5oqISzDS8gQX84opPqtyqXUiKCfGnWXwryVFk8Ug
HGVkbCIL3ydmu5cPDXB328Nif5wJWBiMlu7LJnys/Wb4rHtwNRjMxqxtW6+GOS7u
FOxz3NcIxDhN4I1zKgPJQdOtl3ECouM0TjY/Ph87SsdIn0uHsPATz+mGeUDmjImn
TBCP3rElz+hqB61SEYYj0yqu6PB9hUNUUMo0aOSBNsfSBCrXJOe3QSr+nyQKSydq
0o+G5wJ9ErmPCMrb5YSJpp6PXrNuG5Spvmci9MkW1RCX1K6vDIXFpuwHchxcUr0k
4PFi1/u3wIfeGZ2l9nlJYLUCVWHauujj+unqlVrmhs206Cn7OTyeNwRDHmLEM4xJ
jxKD+Bb06O4njgVz3YtiQHIPiP02GJgnmMevi1fEPbn7DYUMKCBpn9biPrFxkZJy
ziyPQjU9GPC/qpagzd8ExqbIsuQj8myAQWiussb5b/0B1pbk392KAQ7m02V7mgS6
5yiRx6zgiFCz3CLjcwo1NAIsY/C1zQ01M+cKSyVSqsK28sxBimJnFaAghfZmIhdw
+9iFdEyCR09OXQqLCnfbOvtXD8G8/VjmfCWt67GaVAaennuJdHEz0OgWdlf6Xi4V
Q+lkkb/ruDisfYdxYDWmspEpj4Q/KPIK/KO4jBb8iMBep4IXB2BfHMuVU/20JbEC
YWUmjilqWlNJZoTJToE3h3k6WfGmz+2B/rBo/2FFR3tnKK3fAmwLcDMumrB+ASkZ
ymRtGjWVSLELZGoLZ3H3dBVkP09RgmE0tnrmEtWAuBMBuLBfEAS+gUeBVDaxe99+
ya00OBMM0GXtOlzSBaoNTgPNa5ZsWG4y7gc8vRcdcyOtUSuWrRU5wNxW91/3feX/
uzDoOzZ8twmtjRRNTtWSbId9L192vXs/5LXiFJwIyuAGFopP8pHtMkFOUpXj/ahA
1QXliVsS27xt1jXnD7iREmY96f9Z2H3O4FEW7JzMtFmja06ptbNF23IHZ/6FMZ3V
7DqWzNV8ejA+wJLq1juqDsSgvs2DF0oAbh+57yFHDghDYWMvnRjx3pyYIni0ZvKE
7Nyg353ga6OnPM2r8aSmBMuLDsy8WrTy2yM71yU1580HZNIeNrBJKvhkPuZje0IP
lgJurticieP2fPEJCxbLJMeKpgPhfeaKEoBY/SRjPa4HybwS28koyPQE1NSCCCh4
VpRzg8L4GuRo9DUln91t8n5KRTeSboB4+q+2KLksFsy6hDA3jtlVO/1HblmPIGOi
pvhFg2sVFXL7jB8iSmQ0gJ3rFdt3gBQtowlzoGvvohXV3q97swh9djOcFXk/GRfs
zh9F7j+D4rDLM+2dSuKx+iIfebkparqyrJTXK/yTgREGQufib8yrXmqFeTSiTRkz
SxisHlqAwtEzJDmL7LZGShNprIYYgOLf6lsVN+gl82xGuJX3SwCkjuItHdrvC+jx
knHrdZoYj6qdS5zl13uuzgnyZcqOYLSjJVr2GNZ+TdASzpu7AmlHfUQD7m1YzA6W
PUeyMtZEX2306yAKNckvKG5wFtC3gc46ptjjECbLV26WKX1d7MsyCf6kTcq3gN60
di0LUtzgF2/w+cLXPMugoHv0ByGgAWCheCH9B8nCWhdLJx4YZ9HtcuneKMy9/EU5
KZ8JU1jNRZH2HtKgxYMLRLe7TjuW6h8J7B5iXlBfEn8CRhSCFtkub/t1WjhJJh86
GNKNB/UkxqcuWndtdrRr8SrDoRVZ4Mgtghp1cwNaXn8Qwkir+uni7cYbuvgge8+f
E/cnhcfqwHtBF2/HCuKEcvCScBg/UQ4v47PhavPKFaIm9HhfO8n7+VSXfAfpfJZd
hsRbrRUT1rWh/SVmpf41VYCbF5HCyA82Ag7DHviAOJB7X1GKIfP1JRRKuwIBq9hu
Ya1wE74gxchIveUSCIU/ziO5AWJCv+FUFYsCREQyPS43Rp4ULNU/QIrVAtlkwJTK
vqQIB4RBuahqmezzQ2Gh1EAdJnEJOyavHG6ArUKhOYoZ9jULNWRhaaa5PvC/BLP2
u0l6NU8lShHL5NtNHc/SBAYwgImK3ms/lM4YUDOlp095rApEyJP6IOcsdAJUhuOt
1jVfam+BA2TpYZDWJaFc2avZVCkSrBtGgRMrUPDNqW2/Fxuf83fM7cgbQO/bBqzv
ovnPVXVvf0aObqUuaMxNtt5McDZdT1wdAMaUrPcg8N3KKkGgMJnlb/589fwBSYt6
Pg3DCDGQGaKMtAkOdUf+kj8WILyZOTWtwhtD7pZ7gqmMW7Td+xOQkn1HhN2iaKXG
O/wCVUAVxKXyDSuQ0a2fpE7w+k6Cw7Egi6KhiDbHeXe2z1VO7osO04gvmW4vhMbg
ouPDxAzyK+zvuWMBfmvGsxk0Bc4+7xTkQE8XGtRyJqiuBg75SvXS8C5EQgaWyxqC
NMDHc0Y3M8y5x4BGZ0VV07Qix0ltAbyjhivFJ35MjkI4gNfxo3KRKue4UgKlcXDE
rGn7sFjGlNNahXowDRwa7ctYiP5zTOXmfbdI3dlMaQkh+SWUeMO97zNM/iNoWN2P
3fe+Gc1qcAwexIbledG+wdKIoSBI7pgSWkmpWfsdgxcI6ltCuUA8oWBOzfX13USG
byph6BDAxHZHC3mEP+dOX7QSC+vJD5Cpp3itfR7KRFYC9Xcd3ESK925O+fGn15A/
MU25NbEf/jK4J5IuBUe85Rwt1L5Rce2uuzJm66qb869t7AwWhLB+aqzYF1bV5leT
cVTqlnSWgBhKRdCTHz5XDVCtKPjUyg79FP2EXIhJYgLbl0nXVJQocdMzXCaC4z2u
h9q0Uc+uwBcjKluJxBq5D5lquGtClQoKM9emTyEoXkokgbzX6M5l741+XL/hf2qT
N4KZN/BcanCmzm4Sf+fTtEyfn8x9hFnXAkIKlNOAq7Im2FBHNzv9BSGmNeTjZKcw
iG8VhP0QRizad2cBwIsUJpy+z7apMh6SUGbc+R/1MnKTO2nqhzOj4QwqYyCEU9yl
799EjOj4bSsaLHu1tnQryMxCuy5o6UKCdkeHo3rDg4tx1xTYcj89Khpaawx3dSfp
dQb+t68vzyB3348lAlxRXn7u4LUkZ3sw2UjB99qU7XPpYoI3ZxOA781ZBV+H0Rq/
ydD8fgAFxklAR1RJa+Hk9md/a/4I9RhuLF1ZZpzbROAvBHrGf+hf+iiUncnPLiK9
6w07fE7vQMBNYY+gF7L2inY4bPmC3jueoRYr1KhglfBy6/AwnczW9HWbov3HXtyY
QjX1Kzs8ratUxI0rnD/UpRpxM9cp7GCmVBFcohDyhlFzMVPnU+AujxKrrVrLAntc
sV+BoG0huyAUlO9VkM9GXL6vNlkYv2fJi3Fq3AT0AGLDlJp4dFWFIZLMe6NVNQBk
BTaOd2ZYz/sgHxCJ8vDy1JLOJb6L8dWNhq6CnHHdU5+FJiHZ/sAN0WX2s7ISXXYD
KYdzL9QoQ5bvl+Df4ly/LM0OfD86pJUzDLW/5vH2fGejObjOHqfZxLkChJEZpp9S
daNkX5VxPbS6RjBKBZbijr6SRJi5E+fSl2JBaFlrOPE5fpAymiOVKmEsquCbgOOa
LYmoEUndHIsG0K4J1oanEWJcwVZSFvNwpOsvIH/xwz7fUG4EDQZ5o9tNFzh2nMOi
McgQ3HTFOHZ3ePF73mXM3FbAx6hR/6WE40y8L7tB6Aujdo2tJtMtf9z2jy3nsmSD
MsBm0Qz+Tv7VAs+Tp6An71l23EA2XoFM1BZyqtid5TmxodEBWUqGcSXFjXmSTiOH
zGCzJkDe5d7+ZL/p2KwW6f/CvIFIzIr9eZrSTbYVnyCwcHVK3wKxFJp8GwwW8KLn
1yK2UW2ZP+paDPUvJ5wIyerhjHXGAiUbNiPb+W0D5c1Y2RxyoPP/XAOSKnk/EnZm
Xu0QIeTnunApxKd5Vy8Cj03bOAAtaeBY1cOoquypdRWKrMk6CjApN4zgXOQpQdlB
xT6HikthKBKJ81+KOD8nCjI8yBbUHYoC4/FHmLnU7B78pUTPiHjJQ6/33ztBFJ6n
T93iEPQOyTETwgg4LoTm7XaiKyPiRcCri5YBupBWYNlE0aPYt39KtSGBD2HcadOM
nlkPImT/6m/iyqQTJAZ2jNDsEpir79dHi/7EztlouU91feQkGWmCVRGl0CoiRVow
QzMFJRa1xUrFAvpDOfZzXC3QYU0Zs7nmglRqAExuzGWLnN+HOFCdOHEzs0mKpCyP
siGJMf4Rv8q06fiiA4qT9tiOHXwRfYgkRiCI5zKFXzw3SYfDMTxhbEBjKcMVWdkg
c3VucMwo7iOvTOqXBT0hOBFixJTqtEBKGSf6GVnrhi3/ybiF3iCu3RwLqF+CUR27
lt8GWbnbp7hi2NHcf9NGcci4NxS87xcmCvF+Kd1xjYAWqiqpcoLphnBOdwCBMG2c
iMFOA0dGCAvnjheUKtUhg45Z+s5PmUv3a066BPBRUmJIXdyZj+1srNfChyBNFLIt
4rrgGoqsHj8jMIU1v21SgrFfPrbtDBbxhjCOY2NvU0HUmkUEqLundbn4/hL24rWw
F9U6KJSubaiR/N0oVU0NCw7izaBc9huFW+n7QBxolEIsRemjPYUP7xBdFM/EjTj0
ocWBReHWukql5eBpator2PFkwmet8I7FaCmGdSyISYQ9cysU+3IilQzxF32bNfFJ
a2aEXKXcTeNWMIR/+JGNv3jI8y37KQf92bTb5psX02ZZQvFb9DnV/82DzQtx56r6
R+gpEg0h0np53ExZ5/GzwfxSaQu50WqNqCS4Xb37f9jSFPCEnCoTTAYtqi9jSl7k
FubGnDXFX3vxdXWfxTW60vv0YrzVeNIz2rF8G6w2+kQHw4SyXUAabAUpF12JbWGw
QbO9fVlNtAGkY9bmGMcwrj3ZMyM2N5FksnLqO7h/h5du37OOad/4Ek3mVgAX2J2O
UipaLA/575gliqkpGf8ituqWhdwG5RA8US3B1i2qO6L9z7x62gXW3p/pqgK0SHHl
JnvmldfOe6eZuwxhvjLmbn8n289ENsoWFxfG81/GCN0CqbM/WfW8XOhgCQaKYRXy
vqOaVvfR4t4bb3jErDrMaIwxg3i+2Dyl2An21AwOsUeOIYK75PWkhx8FhBd5Y8ts
6QBYJtFHQgdPqbv5zQsVM92qz7GFnjehSrhESdRZOVHoSb9GwUybfOpwDeDqMTxT
EaS1N76KW59vVGBC9+LaM5D2IWwgOvn3FAJ596qAtW5CLtQ8kO3EoIK/1eYv8Bet
rmJ7wQENWP6Yxk1DBRBRg/Pzo3nSSnch/XZ0FYO5Tu9xASttvAk8CVFP3TR0KEuD
/q+diAgTOM956fus/ZCFZExIZ+P98WeNB9ynC/la6HqKWGgLXtTa/7n63+6WUHD9
rCsE34s2uzUK+4Q5+qf/EpVBSqAJoEdjX4aec05epGqc9BEef+YCainZ388k68Qh
HJZMYfTCKGm628EstbrcuatCtPiusZorqb211SPa6I2U9hMd1h0CDE3wWV2cSQrZ
Z2Egdq2rHtNeHj8RqbC3qnkK1RjRaUpehcNOdOY2RIK3On9uL7uO9yTVHBH1c6UF
W46CLLl2c3ywWFcDQ9+ZtIEAR0ALPDxQl8C4MD9FoRkJCvs4YcQDYjNrYNrKgpzQ
FuFk94cLtmmruaNiM8OkEkd+7Zpw4TEUj67Fa62EQw+GY2ACo8WQkmdUC1lb1umj
l3GIp2Xs6mxBTC4uVxujY0cFpFX614wPWA9zB/V005gqcVhuaqabJyg+DMVP6wGn
6+lnuMwO5k+iOvkIarb1VgE4UE4+H1rNodGvhY5vkvHUYExEpx5NVeZqatg/Dd5J
eN+iQqQdwqvu45LT1O3fbGUFcmWA4qq94BPbVXjQ1bwpLuBQS3xMz4fxa8KgLm8o
HRSgmmzhCubHA7QOG6MBAmvI85/nxYgudBHTXpjameNvzfIE4QQpVG4d3Tr8dCQX
sPC3kIfP9EmCcDRSYQafX6vmw+yPGBxSOm5hjxkVKenX7V9FEoKi2/rGVOoaU9iB
+fAMGUmNhZXiFpl9DCFfk3nBBu+9Bs7C9x9qrdIl1XHL1pQ2uaT/9x3Ywbedcioe
oquCxx2TV/ZfPZedDRyIBsxSRuj+j5EdO/rvbw15b3zEHHduhQ37mduew3Q7ebP+
32vwhuDocT7PjAGTd0q473av0/hJqvsIx4EJaWO31gZ4gpSK/+C+Pb19JFjqcSyX
nKBd4Tav36z4sUN2jL69OZlWnPCL+knpcunfubFC90qkIgYtFvIeWGhHoMta8/pk
pWIm3rIequsPbn4U+UaOKVRjaxS7I3XniB7UBw3VHgMtDPvgUExWpfl6e1nqRlH4
16MDfHzGhIoPAHdmGLQue0wSlCoqVl2EakVjP0WWQR56lr3P3Hug+8iXk7v+WlM8
sL+/DcXVo3bPipFWQW0d5X3PfZy2krlY0aGVo6ZM+SUn/bvemFSpMx28k3DoyeIE
Rr7pR555o1T+l32BLuVCNBY9kMhc0ILimw6miOfIHyWhlpgOJYwld3yBEqA47MAu
aU8nnLULKe4QpbSq5lJSE6BG2VQdTUnP5jWXig412U/OoOXHa8CI3lHArsaoTMuz
L3ktH6LyeZNVQ/cTFytsVyj1aqedeSUZiueCVOWpTYJkTxRxff8l+6qbjDzLz119
VHipffYca63gXm53cbxyCzgMsJrhsoekpxZQHr36f4CNHX80UoJqxwcrC3ju5kM+
qJPiR1mQTOCN925bIiBpzJLs74ExcrhzX2f8WDMWCNB4FpS3mVkfhJ8kN+Re3t+B
CJLol8HK7cnjTObIFfPwVgipnfc4wjecUSjrRfelFGuE23/9Ii5m5uu+DITnGqQD
XkbE2LMx78+BBzij25eX5H4aQE5y+CdRxmE96TFVAWVYw/3kbuXZvrNp4Fx9Nb8s
+3bnogueMFSfWHhmtuQXy2hd9hCwZCeStUVDGSRLqPHFclvzj3MlxhVPIWO7TeBw
YUfwHLVLYreNX7hrfAoh+iFyADxJpc/sMNN41z7DwEopaj2BE8F8V68Cxe1cl3O6
c7IvNd5+K7nfQYNLc5MNck+b7iYnM7UXCV+VogA6BXB6p+bfb5YO1LjYEYBTvRC7
u2Kd5nYTSb2FFRCq4DlriMwfN5Dl4pIzSJ1G5DdgAEZfr3zuN3VMA5mf9ydTmgnH
qZMD/yn++55PW3RRTqkN9t68f5hfavBamt9sNuj4BEtwN+Wqr5YCRTKcpfRRiyA7
onvEe7dllySWD9T6gx6bVqPb2UAdzb1SrQZCfxfXtYGWuX90J+VbngGMbFwUexoU
cuY94fXwNoLnG2sl7/vRYOqkcmZ+fwmjSwBeDwDkZhn7hnXUN+DcusIKdCvSNu/k
iKbkW9ENDNr3YPYIpGxDC9krMvp1RVz6M4U7u7QZM4CsEQ8KMQqETp7JDm2fMdNc
7W9kIGnjr4X9KLeUz2E2oP9TL1koJ30Q3q3JS4V34O61dYF12h2NmSUWNymfv3v1
ggJrSWGBil9YYExb3x0yTdy/51HZ59W0fTbdFv0OIkDAQHqI8BK9PKKS25NYFTps
GUE/RADrLYQFisfr7C8d1oLFz9LCTgZXL+rT1ZFFJYm9ejiwc1ahY+UkDRO1evGX
n725u/9opQNPeT7bsfc5IHIHOizOZesnyzfgS9UtsjH9dsM0Y81geZM092dbpuEy
eAvf+Q25SVc2RbhRuAlwnsfRL6dpOlvRcfCl0wuSe678SNS0aLQuwM3a0NN2yp8G
c3FZdFbuO0JngXOSED/f83NUOmGMZT/AfOxQB2vfCxxH0CzHIhZx2n0LBLUvPSQT
CovYffKaggLnkYMrqKJlMn5EhVe1Xg53MEY2JW61U5XPELAMMXPGJGH5IITuc+jZ
9Be2R1Nk+t8VrJWgZdjfInkD8IkQ/5182gLb3a+PyXHnQl27jskzNg7rVN0zMGvg
ZH8RQo+jycBdghnWfpe+C71oHorgDoUZGKOPp0ClXj+RunQI4XpfQSZzPoHm1JKv
VNqYwExcywuAk1Y8fNS804Xaj+iCipOInaD+lGO0qARJLT9AsIFqKjkUYBZEDUGW
SyEXm2SM7bowZAfq8E139LgJwq/tepXxHGARu+sPFew4rGwuNwOQCuPgVI1KZhoq
MX5FYk3l5PxvK9gWT+D9ohRHrckqN6gWMUrXd5uHe17xnXmdO8U1yKz5PN75472Y
vYuR0CxjUbxpykOLEWYmJ7NU6oFW3cpmVq5ch1vOaI56jvhIlR9QTc5RGB1alGcG
Nz130x/dMYQpoI3sCSb08b/TAYKGeZzG3CO7X86tAvcm2lL76s+6kdyzVCtJEr5W
fHpbvAHKd0j5The8RjVUcAaU/Z+5mG+Lcp5ys3lxVW4as7+V+jZzF4+W5YgAmg+b
gHk3pN0/vHNmMOK2r5MmnG3rG+kJ1s0jiNE04oAUVp4+7bcBHulDFeId4o1RPNAr
6LHbnf6EOgTBr5KTXvNJvI/D4wZ/x2CFaa8WFWuZBckm/h5taahv6h9e/PDHj1Tc
KWD/CeSW21+74bJkqNeHgY1CoZPab0HfgO4vW/TUOvmG76MOQaNchJP5BGoN9L/b
+E0/gi3Iaw4dsea7oHaF/Td4qclQMx2mpfCfuvQcVq6rV0arvpKJuarZnuTzork8
+UbbEuKs6/8IANxPFK5Zj14UqRVtIKF5xeXdg4SaX3GvK+fZY/B+j91BBEh8VZ6+
xndWFaOgB1JZRBnsiAAn7rjt+0i+8da0fa2LtaNu1ayTvIJOIfp6AOYjfbxwgslF
onJsVmbpAm2EwV1HcfTULJnQKWi0KA4pxl0ATYnkcRmAh7baLgdnZu1paF1Hrw/t
rV3NZ981D4A9C8i4nrwA0e8WO8LEIWQU+nwTYeW3ZAA1fek/XjaRf/JlXd6RegiD
UfmhGbD4RksYH70JtFeOUNyJuibsJ/t+O22+i2xSHoaZullusVKwa7Zm/TBsCtuN
xi69dj8YQdH2jkAOv5yXqynljvi0oqceMu8vQI+8i2Q3S+c+cGL9qIEvvHmCLr/+
bcHFAWIFAExfjPsKy0r7/Jw/NKTyuXct9zVFf0Uk7yqll71bm3+4cUSMSgbZt47f
ZDvEkzV7FqZpq90MxDAW3b5UBNKZeKdAcHZh15SBG1r6mu0U0QXSQbVTtIaNcI49
tDiOwbLz8w63C6B5g0joJo4hcKo2RpyhqU4zdClok5AgPNLuvVW96QsZiiYw832O
LUSQnAk6uCWMzXggjfX/3kcwC4eglWRceSMFB642Zd/HvsOJYP6EtD2AcsbVJlpm
I7UP2XhMtoeBOcfIBDd6sMhNTXCVSUC6CzqT+mh22vzXi8f2YMTlvRvKt9AgmrEQ
EwTHbAAsUAaJ/IM2DHsqdnLvfNFeu0O/TGZuMRdFUgprvz1x+izCQvAGzFbDZ7lO
q236dyNXaLMoasr1iCed4DLAmvBOQyCGGK2kI5un14dHZV7JDnYox2p54eUuY1Tf
z5rBnHSVOi7ykvgUr9MWVoAHF8EeCA8ufbc8QaW2L3dZjbDr/eJvXxUjMDdzVIrP
9vHwfc0W+OMrC31W6CF17i9QVQcHB6MGQ+QHiZD7Zf7VI9fM3TDQAQn+3hQlSxRI
Jdeltnzov5CxHbUvt02Ra5xHIkBCg1RfL+d0m9HFWMHQnl56+1L1fT1pVOMzrvrS
9ztrfAL6QXwhd5KUBOFlJ+5ST5g7Ca6A3YWeZONcz4QybEl5CMhEygpfpexdmC4v
3K2rzXx7pbyBu5jdKGRpGPRLA3kSHY9wDbpkdqP35Y0fGB3jH+YBjFLh1+EfIvHc
6cpJngcKSH8R6vO8fohnOX2xB7fmGbFS4Ldo2cFRAizTLUPaAkKsa/SNCD2bZTih
jpwBpZgUqYXQtT67ESQMoiXOq8okvPY+nRwDE3BjKT58O80s6znj0lBM4Er/n+sz
5bcAlsk1QRdnrwWYBpxoHrSaGPmRqTbVfZPIycn5dKVAmBgfXQsyiAYXZ9nLCWC3
pWJmXBZFaO6zpWZ51oaJ+WDYy9qhlixADX1ZMxkn1BiRXK+VjoLAHGhbRJvkDsZp
2SzH9/o1iEspIM69kapqLfA1R4DEkkRUPTzmA5fy0+5/vNhZqfUZbAlrHcStq7eD
Uj0qdUkH4qtelXK8jFaLtsxt4mzBNMGQ+9UFUMGNP6/qaJrRRuK01NB8P1INLFas
MJYea2QixGffMAq+uEX9xIcqT0Zm0hZwXXOPL2cd9ccOJcIlgEZ0Xpgl1sbFOfIa
xwt+tI8bMRFIbKa0eFCQhXcHJV+QKyI7TpDWu7yDDC0WfGZoTC/I6aNqyDCi9iAb
e1YLRcDO72ZPLjr8djmg6MX+n3KOHxi2HnANqxhHUDYahBxVptqteVe+wjeU1SPo
YTMkopC4J8L2kBw66P6YgD9N0hH3LKD80tgbGJ7bLcKrU4fTqTfRjeFWEeDzv4QS
izHh2eZmOIHYWBFPfxyLtnew5IiUmnNtPyM+BV9JpWKUOiOjEumh8i0h2HrX2OOq
Yq6LJmRV1GalVDnstwiLJRGKqOWILvT9B9guKMihbU9w2zpojiwZfNLmrvu7BOyb
hZ+Jlt/jQRQ24a+RUpZcgwUbGz9qvEzAC1Ks7M7IUGFvEcRm0vLxdDP2QHmHc5jt
LbxD2kvB6AcKbDoGYi5DZHw2VMmSiZfv/ti+h7GLGc6qISAJGwlJVdVoRflCc6dO
SvS1Vgb6/gSwZz4gJOjR5zYQhJ6pQj8N9v4zf9sTHcaaqY58MaTulctA1b67WdZL
c/cx36s12CFEbTeaaswmSSQ0XxJNy2JfnMX0Crcdz10PAiSQdF36qQkTPfn9Lvl6
smPGS4HyQZXmdLm2vO4oyID5tRh5zE0fyXAOKx2GGZYC3ch9s1zhLjpK5Mkry91T
4mKFsxqafRv0sbdAWVW5lzgc9WzxocNOG4fe9kin1e34nSdtwDJjhP9fOwbfRuPf
z6vNx/4fc7sJu1MeuBxrmnQ7eFDf9xvdQ8Y5Fx62ayF0obQB9y72dXumuFLP2Q++
1qybZtTHCPrVNiioigpfQ1u7L5dnS/Wa7Y7c/4dE3QGRwT8/DkQUpfs7QVa84Kq9
F4DTpzMH9Og8C0Y9P6iNEe5SgDfGdg78s65ZwEktDcJwBeNs2tIecuzeKS8mqn/8
w5ZLqcBU+P97Kl2BO/hNi77JhCVLr2cRhUqq5Caqn8rOnKR/jQ1rZXL2JGqUfxDg
eKIru2zbYt3ytZwFvvNCiLyeRHN9tHD2DEy+1S0uSruya0HODDm//QV81LZkqiiR
dj3MFkMzpafuYSTESpa2CPJ9WfpJzqPerHLUqEwcxvYs2SgXt1ZqZDE/4+o4WUn/
bBCRLsqFvRQXtuUwqdOyzPr5sLa0dHhZzVgliIJ2QoML1Ft0K3iN/hby35OqsGFc
XIu8TbEFMkXb9N901AUM927oFGXsaYu6nsd1WE7UveGOWqUPV8abtBbvmD9LDKM1
kdqcHGdXy7ikky6udnm6z48yFpt4a5zf4sLM7r+n161IAUu2FfeDbM8FGYSpxel7
3SqbwylIUZY/uBdjE/yaIc8ikYhtz7R2ruW/dCxhj7LmZdaAAhX3Uildc8ScQmBh
QjFo1R5cxs78tkzTTm7REvTbCxU4AXfdds9pB+nIH1YocL8FG7YxGEmRKaWZsVUO
h16z7+ZpoGuw9FJhmSvcoibJjG9BhgDjesvmZJmDzk0ZWEiOGi9QHQdrGycblYD3
f+1Yx1tmpnZP+qKDVb3T+weD6KpZn+LirZTbasE05VnQjru0bme6QTzfeQTGXj8T
IiLfx5ABeR8BLiJ0GLA8b/nat+jktvDJO1wt26vqLPi5+Mgg/3iVTuo0PYbgzc/D
olDHpEE8MNedICvSTYqWogEuzKHNw7sand7g+nGfeIQKYHU9Zk7zvRYnKORlH+vH
iqTuWhcCLL0q0iQszhmHUGa/qctusWHMW4NVTSn0rtXehfuH8zz8kmDPEAZIatat
0B2VoYF1GuGgcYRvnSisCDUo1Fd0l+pDDnMFKVGa+FAAFHyQyDxXUQwQAZZXaOtT
XOFIDynoLXVw+bL6oefC0rVr8GpQpvqtklwyJpHqG6YdLvbCpx3XQigZb3lHFK9T
IjM7W0lv4B3BpL1nXCLBWo4j2o51bMUsK/ONNfB7rO6DiC86x2h583Ka3WDdH1EG
X+6kwWG6B3CMxPpDE+0osytAIDeS6DoTpegws3uvgJ1ZKOtYllGgis7wS7mzSF+l
G1aKf9nD3A4T2pjAGBZe0GMM0Gl8arzHv4e2PqtEmjkKddOipPt3t0YXLqs7PeXv
cLEyhEhdIhthyCX/Lqg9Oe+pGHIYOiFD3qLnMqC4+y20ifdL98nmjmMMzepet40u
G8fdLCo2SaYvJ9ACEZJU5teCZ829AWsbcuUNd3y24iuHDtd/AVBn7E+yKs4aKPxz
2fsMF+JDjo1LjYTA1Q+zQ/FNSS8xIHzSO/AN/PPDs27SEwaRc2fUjITNtfAIe+FF
yhbMhA2t/b59QIEbKYg1oK50q8TzHVyQao6xXX7syAy3xV6gH7g6FGGxM/hMlM11
j7QbuTYJZCd5+vauDwXkVG0f9b4qnmhFuUg6cfCV4WdOXPxkDmXAdTV0TvIsWDwX
BYVl3qru5XFMfik/B6SYIjcheRFy1ja0xTAq3ZqkJO/VFDksLWiZjA9iv2jlVQZF
dYXV3IdFmdGAiGJG45k1H4ddLM5FqcqpKEnb3fMuhIBE4KF6wWs+q8CMgz+HyHQA
VPKAlgAYKyfLlUuuL3/QzYNzUzZtvZcl0Vfl3Q3/X0We6yWp439Lu1Ppe+lupG0t
7uuzPje+QOVv84/z4wIC7v1Pr/Igs1Fx/fq1DnrTIY6HqONc8sSxPj/UWfshTpVK
juzoAew+xeHf/kHQKxYYjReWEXrhl42eZnrOBCH8Gf4Um7jtK0/CBffH8KJFXIYA
osIL9lgVf8A9HvnbryNX5V2Z6Y+WkXdLCTm0Lq+Uy0oKj8dVLRqGNh8+6xjRLW19
dguZ/vIMk6qxRNVIRtJE9jckJIlUwfLeZTu7FA/SpUAShj7xgHHTXYHRMvvxNxvw
c5RVAu+QbU6MHr/W7Iyz2VJbujYOaHZSIWjGlTaYyX0P2YUb7Da+BMV0crvEedkB
Sf+DpiE4aplPIwVngXVZlwYqN0yjumQ8j277Knkg1KAEPYKypDvNEFEt1LyWrl7/
HSbAkzXqPd6i6561ujucNIowLRnNbDzCMvC9PPzOUlc5PXp/yL8gLiOfMU6txvpg
0skFRQRFegQJOa9j56FWjHJwkvbJLVYG3uGad7/pKz+dNN32+rwkziSkK4eoPwPp
9A3ioGNlcgmpYpHimeZY6tmAKs10vJra/SJPGNIkCteba9H0XZd/l/tscLTJXuKF
Tkr004ZlSouyXayKfOmkbQkGCnvHm9z08UYBKfPWy8Z6hvRpwTzetjjpBdOVfvNw
d6Wbe7U1cobFa9c3vjE8jKgad+OKG39cVyCfz9WxMGwY7YrlvYY1nFbJgKalYdwU
RnMo1V39QbOv4/CsqkmdobhQzg0CqVFNJLEBDg5qsyKuy11zQVu1hP0iRr0SuXsy
ExvmVWhz6m3X6Yze2CsGP5BsSG7c+uXucuC0CPzke8AVRJ93mWrg+aV+CO4d4Am2
ZsGu6/Rhk8cR1/4duPLDc3eDervXSJ9dIfJKWVbb11ygSjh6Pvcqmca43Pgd67gJ
+vZOwCWcI8H+LU1Qxq2DDrNXqeYStsXrDfTe52Z/lxvDAye2Bt1zJtX+QcKCI9XL
8fv5iPV9zNJ1KBfgrOMCt8094KWjk8cOjOs0oYNc4Uqyqfww06wgBTZlX7ChoguK
xrINr8rWGm4QpS2buYyNPYTw8IhnQxhkK2SwqLK3A/U5hzbyfWY9VlrfT4c1Zk7+
dafDfgkJoq1FpfS/yt60ocuHhVpDo9DW1RReJFqQLz9HvD/eFYTSYti9bDrpojP7
/rxf3gO57UYB06CVQ3UCgYQ5xVK8NoGk7MABAcyCGXqZaZumZ4MlW65BKo7JNGIn
K2lxDFDLaXLZbMJj12wVCj0ymGUadzv0UXM9ABGAromCuEc/3ePChXHMGeFuDPIF
inI2QqORNLlba6SuTd1qLANHS8M4uY6jIFpUxPQpR7ZVr/4BZa0JWZljJMx+GH+r
qy+zxmcQB20xX2wDr62z80CRIcxKtXUIvni/Hyx0q1Bxy5x+piaDmikb9VozwmC5
lrPDly1+9guBYrsR8ENY3VZXXY/Spba96Bf31law6UtzjyhH2jICq+0WCW+AarQW
+q5d6Cu2jDIOa8rItbpqFZ9EMejBoDLKc8rFtyuAs0b1RzLF8VTG0p1VixB5HNKB
iRYmbU3iStzh5kQCFDhlI4TVG4lbWWSibaJD6VsvB608Xzuzq5HQyVwIFCS/E8K9
WrQ2bvN2ZBVTj+jN9gxFrR+v/TOc2sS3zQAPR6AKHIUJxolnVk8bJ+qNx++oyd+z
NxH2woNZFwHD+J34ySBa9UVYV09K963HrM0KHGzZE9zI3NjXJPPOhmJmz77e8siu
+VxSrgAPuxoPXbyC8Zd/zdbfFjyLt4jfS0AqMxMobWLgdB9d8Qsu68EmxnLfbyNP
KBJHS4eIIAdUI+ZScswkJisi2WJbqsvuQ/27WOknL7GyKoBCk37q9a2I/dTunOaA
oqHy9XxlKVJhKjGVR0YOPnmcnNFsJAiPTLcpPWjOIHxBL0D5okfF4CmYDrwgfIS5
0fGKEfbVli3lh5yHClM6A8fbb1D+j4bF4j6rR3Dx8+NnUdGnHkkt4ij9UHrg3Zyj
W4ymNLtbdT3vWagulTA1Avii+yOHRmIEDclKUAOZRvb1NbSdBDmVlTul4AVVuV/p
9AxJCbPl++dEt75MKYzxjGr9in/kSZ/oGbADmmFp1mhjJ6vj1sxZYzVTxXb3QhUs
2by6dTwEhVKDoBCiyLxei02fSWdHW2kuEXSEGv8KlpbioGWpo1GGFWnuUVa2lovV
jS2WEqMWSTiYhf5UrZqBCt4dEAZe7tuvcwMP6k02XtQThT2jtLHP+3kL6+Xp49NH
07Op11wt6rZDZJvtTUvxyILp5R5yi+jBv3sjIegiULOaEhhK2eVPw0owaJFIEQLS
CdHMkO+sE4gQ32md9jQb+3Dx7zZ4C1qeonH8+S8QkkC5YKW6g3ZTJ77BwEIwwsf5
NcBunf/qar/ETC1+Vfq12Khn4qBpZMLOusEo6McS8nd7nhijElk1Reur+svuNbIL
OiKPExnoBYPmjwRCQxQityDxktIwb/AmXpPMy9qaKyhBEhEJyrD8Lx1Ofzebqym3
+bCzOLxCkThgcuEDyog09QtprfqZ9/Tqcc25i/7+4KYL95kqjlmcnz2qtxK9TaKG
KRxyop/C5J25uftZtQKh0IVla00L8fMIhCR47oPbjW0XdZwYQ8QA28cDv8Lf0Pqj
nPNCAtpKC1dLP5zCedz5PNfxSnv2MV9QKLFR5jlFBkSlIrxbV55UEgLa+KUF7plS
G9Yyey7K8b19mGuqgQeXkWCyUV+awa0CcRLt6562aZ3aB5lqnH4+qKb+vTz9N9Ke
QmKZ94rVL6CK568YD897+iOO/0vKqUOOyjFaPAEUhbIbHeokVePNMc6dOYb7K3Ho
hMd0PSeZ78Yq/UokvoUjJDsWEa5KqxmfyGCAFhItS1L2kPuhi+XPy6yntOk6tiKX
snqgNMT2YMDMCgqRj2QMbjqHL3EFPZOIh4g0nGy6OSyGtFIFG4vpxLTwfrjC0nmT
sAD9cEDfilXohRwXNgo0a6cWHjK/rRMakwL2Bdk+hhNoVTLNY/YWdqsmXzAtIfQM
aRuyyHQVqgV0MT/Z2MwimkRUd5010RayWUED2or33kOnODUAyHRPbvE6DvLskMhz
tABmodhmHYEzHdSvvGI88QHyQWAcrjZ8BoRj5WzgtdF2R/drEWTUqyYUnbb7TeTo
+vYjRcQJg3m0Ej2PDE8vT1FYvf3CurKoCGAsBEVYuY93qaSN1Et8uudJEVTrE2aa
GBIcP4v2Vj7k0krPo0JbWbrnbqbq0f6m7rdLJVRHq1rDNwO0oLnSLBOwpEkzDreA
xGbNQxNQhoVSjZfvUrqlkQNjNbdBjwlyNBw0co6JLgbdSCsa9Pko3L+TPrTYAyns
QJseN5KkdPYrSv2dUinU0Mu+w9XJ/udt+OEuRHUb2kv8jkQWX9AFzTEmP3fi0twP
JO2nzQwi848jmKQo+3vyhuAfuojYEY8TNnr+aqQZ8CHDj2Am6Pff+rHY9PRtiG4Q
fQIzAwVP874pwAHDXzwRwhp6LLjGsmShAj9sPLaibg8kyjgve1KBeomEAwcEyir6
0bzZbeQzD3Ab1b8QA4ajybsf9g6g47IxIHA+6ST8lXeRQMkTwVyzcpxB0KPMx59y
2UoXVlr1fXidK9UYk9J5+kmyWgCDI6jUw01DltufTvqhtLUAZWmvTDIwIUTxuBHV
OrckSvGmnv1edxPBx1TJD6myzg2vXQOOJBq2cGDLyK6CviuXekUy6gBUwa6hVdpW
Xtc+hF1PWjoxfw8HYEQCYndVOWqK7NZPAILaiVBvvulmDKvvumkPCpaDzfTJbw5f
BfTw/mawl+3/j/KQ+/TLqG4daP0PcJXqmah5SR12j29S0Mgk8YsS0h538FGHdjHq
F6frJarT9lzgdA8cxsdgn2NcddRLiwohPj3WcMM80RVWDzWattxQHV5JYUzr6dJm
9O7lHrRpFMmzVAWua1DeYTFe2sw8cVqkkL2uvPrd86TNRRjN/f9zQXU3cQaxm39k
KDgoYxsnZDs2LEIW4jGZvGQWCFvn65eAH3U/AsHJ9oyRpyuMoDj247ijW+snpb3x
/NfrqgI+WgAB0ccNSC+cC+kFYibPAaj3Ywudcu0hs2SVXD8vNmbqqVHk9Q8ByrD8
W4IqQgaAgpGwY/d43lxFbxdELmMrCQ5k547IBmU/4FFdZ2QfZDYjZBtpAz5q5Ohg
EBeLHjgY+95Oxq/e9umg52COsImUv0ZG1TexDMwhQr2aX94ULeV+QgJUSZkK78In
iji3Qw9xhY61AucGxZ5ck9gPiQQb5+UaCMZ5M8Q545A2c8RMM313cpA3t5u9phmf
Z+uZVDL/aWbPctixgXUJoDELUYwFB2uSW5F5U6SHuFngcl1KKumopsJozOdmbgcT
UnVEiqdzPOQ86B8rCALpmYFYoOqrekX7Ye7BrKuSwh3hRZXJWVHWrUUKjgx2nTd2
gv3ypd7jnQu3GdsGmZaDE8CuY80ObhJSVorn5sebPOXtTB+6PVHUvWhh5wnlqu1t
eJX7hY6dMfobOxMzhE4j38tlxJ93RI4TelXgfXVKfqsa3CUAMD4o1AeMhnIDBaT+
VZIlZnm0G9VmCsiala9AHPH1PYH4WMuvJEOXzZozReVGMkSlpw6+f1oRGYzF1o64
YT/FK/OdjqHw9LUYf9dvIbMTCWtwQ5mSHkd/4zoG/6BJQNTx8DXx1evYsuQsUNm6
0YlwIwebxgwzxe/N0ugc2oGPmGycQuwlfRCk9q0te3FmF+IC0vUdfJkDy4RcFGCW
jTR37BMzpPwM1WfdrTH54Um5GlAJSK9N3jIN0rzlpFP/BZcjj6azAdJLXjl+vh6m
UfjXt9h7/q9+SraVmqywrgIIJUYRK0YHh6EI+qqBfXlRDKzNEzdfwCI9w2ucYJYS
46+N0QwfrC24OQDtlqXnR085D/KVOpEE+HfAL7MINQOjYFOsC82T4GY1eGCKEWyb
58w4X4huV7AWfT0SCMwQBnrTb5lLER9ytn60+DXbZad9zZReQN9PrabrozYk8jrT
H2VPVqI3Qel5S5qVZSe7RJssWuwLeQ0YUHKFL0j4AV0LSf7XABTf86ryw0WfECPe
yAUgVHh+HZqgSVdynEUaFQNZOgmGh+gHFGqZc/IALAYDC32ZqCVqEbEN+LeC/XhP
7wBFYNP+JInr286Ymz7Tz1oVx+8L3cd8zUeyca13BwsIrcE6KDO6gBgXHNvuENCT
GX2xb+qq7ln7lZtoIMk4rHjyQAVYbhXgZgMkv9hy40wDe2AyHflxDvtfiZ2YGr9w
w5CipNp9jDljdpZEuSWeqrXbBmlW7HX33idkC9WV08tVfvySm2Wp8iWCZWFv1MT+
8L8tbKr0IkQUaexc3TWGRVUXHG9rcEZHm3+dBw/XkMpgIptuuYrc/vnaxdxmSTS7
Cqfl7NvZarq1lqT5OPt4PEqg1E6dJ0Aqd70ZEvDJkm7U/tPq3Ap74V6X37VLrMBw
1PDyQs/FdDEde6uRYOa+FvjwT4wfeRhEIfZ5PJeAsaXO6yUl7Rbk7CzVvju6ocj5
GgCA8RsHmZxRrBPkR7rcL1pTAA+8xD3uX8xBAS7EiS8AfrhN0d69q1TMrnD+v2Z7
ot14gZ2aKHSzV/WbY9qfr/I4wdAfyNi2GCcgkoNnz5JSqZjtmOTjp9w5V8az38K8
Jr2PuZ2Kh79UStadWbTSFK7shjbs5YHM4IckZOzLfMQR92PXUxaxhhh6sYcV5M7X
1GhSTdXNQ8tnNg7/Yd8RrYiGt9r+/Dohz/ntjeSaumUrrSPCpabzJEvFf28DxlEY
aOQNViHUjbSpYFs42lxQEfQVJRUVkUZ/LSMzAJJXeMHjlpxeo/A21SzgU7CnCAv+
oHwpqfyhUOPUXjlFg2/4xiA9SQAtHComI8NNN4pDCAajAZ5dI0xZZsn5a5PMMYx3
0wV4s/M+MlhwxXhsPxcsrGMX9QtNTkXZrENEIs5vIuoGKCjFB4o///87ijBPr7W1
NresytyIMNcqIR7JSXF8/xxCPJhy4Bw7KD/BNjcAwnNWvBpv4B//ojJvQY9BhPit
a4q7+lydJNlfS+0BHnkDm5qc/ItyTRGljm1dMtd4rOMec7L/yJ8CRKmEpyzrdOY4
84nFU2WQ6yZorZeV/N92/0m1J32JMwaBTokYUZV5pGYRgg6UJTgAzGDduzifB88N
ZJrOplwrLrPUdAFdAiJNM8CAufWZgo/oAwFFf2xV6mj7jabqama36dA/JZa5CJcd
rowdcyRScP87GOxNsMGB9II5PlYD7CYr/hyFm8O9sMG9K6W4QNn6IORHqiAuyW2v
u4G/xkDT+LhytwvqrNvYc5Km4HZDA2qLNi30L38TzTcw7UInnyQvDxU6XHpOlSnd
Y28MqudRAlkdzd4sZnianwcYm4C+Y/539URQ7ftvr+r2v6VZ8yDdpjyzURX4+EKT
ROJUiv3Lie7kSd8Dtbp6gWUrHv3QyKqpIVbJIJWKllQpv4uYXMWMeQhaLYbvTtiE
StdOeljC1VjSTmn6lEzEfUjDBLP/prD+hiHOQq+XmVvYZmkRc2+3Mwh9uRuMAFch
KHxYpZiN9j5itei5aIBHdzv0l0KtRYaKFWM7phDEPRPXgOEPwNhPUkm22Dm90UBl
1Q8m0zer5yxUskm26tcZJJadGS2vW/DGEQvlV/YfSolywV9zZ9lGp/ZdR6SrAv6w
49xyJnL/pp+fo1acuZOIOPozoQuH5g8NdcZZcSP2OCflTjJoJGP0gj352C78RyTw
kACBEye74xpNcE3vHm+oBzWcmZK6BJJgnoJy9i75b7bvMALDvQBwyk0gCaz2g5Ci
IjhgKDl4MMIT4JDBptpTLRE/0aZ5W3uBmx0TypDVtcW9PtdB+hkrwHZnlIkvXi/1
Z2oDWhDdCqRlxIt0nezMG/A3w2Nx0QQ4WiFs0GhAkdqtbDe7e0KhXBzDGSbTq2gh
KHDm6ZcpspKPE3NWvJzGw6Gsy6cXjuQUVNP7+m6MrAH/5/oAvoAaex0Fe1LO0tVT
oc+eYsbpErAvcaYzWskEu5NNzzhg1WX7R7cVyK22ty0i7HaPXOSgDRwvfw1P3rNi
nEBeeDPSAUGq+rnU+cZo//uDkly2mxnmDF7Bw12dwINsGFFrcggsCKxEd5IWhFEJ
uoCb5y+Wy/j6tKEj1EWqcuVPg4SDfsmGlbPvG+FaV9vFiqs2Nxf6STXxyMj6+hab
EmLfFdOfQ0BnSUEOL2U60m5zBcEG3ocrhs5kxRz6q+tt9+eNBVzaVXaa15Q9GE7G
BNKv2Duoi6VeFbo+gmAsKJsvOilcd8KlFmvFeiAwZSeIE0qgY/ZOdW9bO4oZgjdG
j/8fEgv/d49Eg2FsSfJJAcTYIo0yN2XdcFOE0HWVI6U3h/uQ2NhgevYISxHPcrjO
obwWiY678Ov0rDVgixtfgqDr4wDIFSaUj6jIqc6wu35WoTEnteVdSZO/pCy1NtsO
9GhE7BYVitiN3RtPzKjmhYIhqcanH00Jh3z1jfWWBsqrRT4PZFEMFxEQofQzZerK
llT3I4nrcTrP4R7njz4YfeQ6R3hEgfqVXeJfYIWjmfE7OF6InY2FNYLbsY/FpHog
9gidipp2QElaJLMk+q83mi0j+K4ZqUtlbCgQEvHdhrNBz/26ab3F2lsEvNDW6DNh
jjuzcwCzVSdjrBIi7+ABcKJQiVZUIDJvey/1XGRx1CRAGmES68wNfHMcT98r0EhY
907fM4Ze38qSaxP/vuBv7Jl9o+wibuQzXyiKdjtwR1X0ISkyq6aRROlNnMIUBVbt
5M1uPrfUkfAF8GwFxAcIUXxOt8ElTsFV2RIJJihA5t111izPXBG582jajuyn0V7n
4eQ7RRzvY2YWWAPAxGaYHm9ngUlNvAue9b9F8Jn9U+EfE1kPC2sBFeXw896M8Plo
Y7/UrlITBhD+dLnE+PA9rvH9GGI1yHRTRyHn4jSPD9yaybGk0WGEHA/O1SCxaA3h
Le5WasY+28x1IWV7cQ4CDCDblnq0uyKmo4HMvAT+rueQ0vvqmODxyYyFG8HHFUgO
beFiHYahK+upLwjsu/3p7L07Hnk68YkJs8J4MTU5XgBmWijVaF4igeVIipsCvOOC
TmjHwR6TR7C7EaqtnFq/eCEbshksilTiDPLn1f0YNGlWGcBwLb+FFzYp7Q9L3Ltp
iSoz1T9lDuQ77J38SA6oFiV3nnS/tqkeO02enNgjS/+x1ORiGmUo/WI3W9JITDcO
lWY3seWUfZqHDB1k617La8hDxr4PM6natpsn8LxHodxVme43azvh2vUnoPm4kbL7
IT9XZjW+DKhFDUb/fa5+yBE3gisYKgAzjydhZwWF2g2nb9HLUo11sJPZuBOSrrfI
LlbMD4wR+/rMIfnkgx0W8bqmn5ILuNuem4OE1BTBFylzJ8FLsxWQ4uiG3cq9WkEu
Kpjpy413UKV0tNFB9lT+dN/BKypoQ4ld7eAXTRzySFgHk0iYAxeboqCBHKmAi/fN
+lnKNj0laJoPfNeCYxcqz3tb4t8ABQ56TrWh8058IFxr0lWz0bsdKarNGTWGYvDR
xw7IwosrRhmaF9nUDYmVppx4sy5L6Kt3Wti+fep5nUdH56Reti5iBYRm5NuNXjFB
jrseXf5K9LCRrPjRVZJblLDAn16L5R1fVsRZ8erZggBJ4GrvM1i//11khF9VnKQS
WzJVRUzYKqim6SRharRY491PBKQP0KkBxARfKjhfneW1ee/CqxTU3rZS41e6rtSd
s3mZL8G5LIvcm0ZXQXR36FIpQj9FASnitpKp5Qr861RgV5Hs28/OcjKYHCzgwS1d
2bgnW2jtK9h+FJvuRZuvur8T2BlqnxkpGikSKAylEIVTGgDWq0Rhn/NN44raenKS
VTFzlVRvbA3kD+qPLa0dxIdxaXBOQ6/2Kggt5MD6rIYNu20Htrb6hXeE4/CV3K31
ZaykYF5kyE7LXk1eN4SAB3MdbDoyWfk0hdSCrKSNuRHWrzNjbOyLm0EZe5UHjCz7
T09Bf8plzFXgs5NVSN/6ds71IcPznWNicM7gL2hDY/Os5fXbGc0rzqU8nqUTcko6
BT8GDiFzbx4J2GTCWNOFpta9biFbvEhbEq2RT5JqU83F8FQ9P4eyc1nwmfEMMuJo
r0iwd9PlxMI1sUmmSOa7k6/p5/5bStjRBumweSBZ8+kSi5WX8EUb27CG3ARF8G9i
2J2X7b5qT5jpt4KJ8IEajp+iv903iN0jksi3Rw33Gc5G3WjTIdM9Lk/IXc+kYvR6
R3Pr2B7xBpUXAO+o92LdNlTWvrTmD8esc2KZnTa9E5hkpjV/pq4T8N/OetK8HYva
FC3OFbSN3iWBexYJNdClkSoLJyg2kKX5pS8iWqTVnuuBtAB4P0JKxXMxITVeNh47
dmaUPMLsEIFoFCY/0bihrzfdBEPgk5ke7F3qj8Tlx8HPZPIlr5KV8yruVo3wBn0K
RrShULrP1zAiJ5HQ0oHEuW7cQvsYuekB3ISqN+heJI8MR/KXVLjVYOZpq+XkvC/e
9dUMdeDYzHEgMiF/JVieV5RZBaP7OlWoj9h8Vnvc11tnH7Gt4I6xQbn+oAN6LEAF
nhMSgHY1+sYgXRJu72/QpKn29/x9EPabPY+iqM3+NgrShMmUpGS47rOvBlBO/Iho
lg/az9WbVsKdTgfmdAjap1Mf7gj+r8IQvoucAQSOWqRuXkO0MbpXngZqOz5tOfiC
8R4U0fO03trBaJveFYGXdG6LG7ahwg2KdnkStk4Cp5HAIm0jTYLbBZ/l45LK3S9H
/XzT4e/xXKP3zpBgsXdTGEARLBXVAB1wicH7nzp6wpFnEfz+cos9pbe5wrUlxHXd
i46isvGNpRYYfwfO+mmU/NFvT7V1li3t8qEfdSS3pQ1rmI6DKqELHtKWSVutnzUy
SsFgQx723rBSX2IPzpLXKZzXVSwEN4nt6x17C219hPN/Rdgzcyw6S9+g24MLWNvb
9xg7mdQL0O97XNTtaS8yPg/PchUpMZ4fT1tMD7SEAT/yYbL55RgnUdazyw7lS90g
1DaMBeJqPKB6gf+ZyYnEJsC1+d5Fh8JQa6e7X5pdcMbuKWeNXmxrqey8i/NIVVm3
En4Gq1YkLolIV9gHqrP7L9UUSmbX4ogg3/nRUdZZ+dc5X3sJu+GeQAMfKsBoDwaG
5nxf8JbysTqMyr7hI4V2FwLF3SPPsH4Efq+ny8te19+WZqi2nCeRN2ejztfd6zQn
+uNBiSjpldxYcFROa1JFMoSEyqQ9Q4wHCenCi9hxgCn9NNRUjL5uZo8S9BSyaO1s
bxT2uA+xSPi3UaZ3CV+3ZwPKvfnHvImqZxjL/L8Fvrpts8k2CKMr+LeJ0iJ/cMn7
8C8/SNpkMTD7z1cbKOc2ddJlCD9nWfZfTaPqlnxW/RHZpEnfa+6eh4w3Z6b34TFb
twK9iEHW6cUqxHmvYqCt6laubYRfEZc9i80HmRF3nv63T3xbIJty0XTkn4RZUm7E
fng+vAXerau6O3IOJbo3T4R3xfTxyMyJciSb7mEBNmfuky3IEvo0z697OUH8doLF
EmksNsUJkd4BSKAVnMfqfk7Pf0Fi27MOgvuPbLyjJRg63Rea5jTTLDAepuwkP2IK
cEFirglCk1jCZKjm1R8EGrvbJEr+tC7GbawqSdLnwQEstLTnxI7cRBcUE9yDBnr2
tX/TbcAKWtmCl8NdMkRr2z+OOiDrk4vOIfQ7b759Sgb9CpR5UKZyIcRw/1UNFVwz
3gi3609BlVPyslBaqVK8da4BOfgqBWIvJ8tcEt+5tF2wtCuFuW2QpSfGq1Kbjbwi
ttTgkvCyA9lKkrQ5FDwpZMhZW5btLT2P9tlDRJJ+kQuD1Q/1QulfEWC6ueE9jQ9U
bAg1cx3QL2SbA3ZHr2GGgCOWP//wB3/4M39bsyTHwMH9zM28KXlR3sprX4bP3nVe
4kIUJWjYCoqUPyuXxThTF6BLg9jySG5G0hIBJK40at+EHNuaOyrKWnqvYXFCiJki
AB8d/Z3gIZPwXbPftvlEzCCzOzEpp53DqA8exJlwcMWyT+9NwNC8bYNqiwBqwd1M
4/Ua3sHJkSn+eXvTomFcr4rEj3EN569+9+VsruJpPGiec1P2FdUBBYmRdxIzD7VP
zVmLpxj2SsqrdCOSF9RDvqaLw06Vm+MGhBoTcc5lY9JkCAz6uW/wr47haPcYUKhC
YkBSkINqHsJA6epev9iMd68vj+fC3ZIlEFcftgcRZTgu7JIy8rpIFebMYrKiQbLG
5BKVXF4F9flSMrp8CpxbAiWHaaNd10KgRVSUfT2KRknX2TenEqDlgvcx1pZNa2e9
IVC1LzxJ7wrJ6kk/UxRNpQdc+qIrtv2Yw8yRpmc+sb+ZZo37NVRgBMBL6Ydt1aHc
XF38ISW+GYF84VBylkQONYU1ylV1NM/1D3aD99GS35MMG0iEzg1jCAdVap1YJFh2
7TXkxcXBRl+MdqnyGcZOYbggtPBvzxjSTUOTvgWifQC8IKW+zqOHpxahjL0j+nF6
yH4pKMQ53F1rTPu3ke0ZlG7kwVrjf94q+auWLtFKma5Ct4nEc3+02LyEspkHWjgj
d3XQ0sSAp4VcHxB0fwpy78YhzM2EAe3RtGr/08VLgHl4AJY36pofeyo5T/9Mr7tm
A5YY0imhQL/4LRjERQWkgHGdZZOBqL2S/zQLfjOacQpTl6rdPZDyfdkTI7buMXD/
t1FNr9MriUgASI1ALKhMvIqPur8gW0FUGtCHmbKha1sl3M+c0szYbdbpX2awacaP
ZIvYEaS3B0S8C/q30np0q/Ejybi5qqYvALoUTS6BDV3NP4l1HKtxoYAkalB18QeY
MEqS65a6/Ke/CaokQQ6Km+4W76xDW48Ml5udzvLYxbIIb9ho5KlN1unEmOrAaPyb
ok/Sgdbgj8gWp4VSfc3v8bMlT3cDHiX0zPuGAFxZiYp+/6q+A9eLh4DK6HB2oA2t
KPQOO0kP9yzK4b5U3VVJW7FUV/I/EQ79T4r38tUeslP1gDjQ7bh3Vz1/hOZa+YM0
7ELk+GXjHJEUlPEuogvbrB6pu6RzHhPfEdwxf1bKpqReD7/srUOGK4TzjV058/+C
bhgqKuJmKVD1P3djq1hXRA2RnZ6rChjWbBX4QAJagFCK7qtjpW1+k4IDmMzS+MhX
7o4e8mNWjXvkMqHWxBmt/gDJ6Awx2KR6uDkotjUhwUZq+jS7fvXlyf3JKG1qyulR
MOota5zPwGvaJhih81dTr9tB46G2UtwovojkTyv5D9VeY9HLAhPFZ4LiYueztNh2
hKevQ+7JNbMZXKQ9cMylaCAioU+1qG9iAOK+uiYhdTbOAPtkLxpx8Qb9Tk0OgXbe
3wlZyYLluob258xqY4MJsB50Nfro6uikLJNOE8P+LctZC849cymZBIVgK+0/7ren
WCrfQ9YWna457aK1pYpDxxUsn0FVc17zc+8scuiOOmcIe8yGjysqT782KFf9X9Iw
OWpTP7+x2z1MMxgs5MuNJaKJhbH+p0xJDhGIccLa8DmtJiHZKtzu59BzQrW60rgT
WfLdVgPn9pqQeKHFD4UXIWG2d0T5kIXD3AwbzwcueUUmjcas97mD7263o7ibAxwX
DjaZ+94yuo8y3bXJRZuc2v8IpWGkRJzXM84aJ/tUGQCpXUUBaNOFIBarw2wTnsCq
c16QWtHKMKZZZsho+3IincBxOfH9a4rB3IMcNMBXCb46EBbbr8PzB1ORFUIW1Lq1
x0GDusZSNfPyexWwzIJtpvfWukR0xvM9JdFB5yS1u1KjX/0O4sxdaHtd/ClRTx8G
We+7ApYDBhQG+/bHf4PvVWWEMNkCPsVQNvs3TbgpS6C6aB88mqN6mnt/gGV2Uktm
xWjar/PjtCuPXGBzZbIOrtllWasB3ynyxntnQeWuyxhB5x771qfqpHlUZbZlO72S
apgxs4S4gDF3bGs1MJymdYHbRsaST+iPkRmqN0ivYJlFLgr1ajl63M4eZ582PbQD
pNLv2Mvj4EQGwpGiNBtU0o1NbTxrfCVaeMKI5ToIvq1JWTM4rT0K/yoBsZVNPyTw
sgF0KIkZM3HwpEz/AHaWdBGhzEyUx06PVn0aODRs95bZo1lmUWQApuaxPqHlx0T7
rojWob6XR8iQr2+fuCsJnHxMbeDb/Ffc5XRNLLJ2PS2OtoG9kci9ocq4yZ3rNF8i
OpmQI4nRuy4ceGBE0xXpZu7h98blvCrtcZshhOKOJWt8e1/Nrbc7cQyFtSsjyTQO
xa29ZsI6MMqaorzgj+1Q4IzfrgbD6756sBrJC5pX/l5bWP2X1guW3GFDPVbW5pnb
ik5Tm4eik3BQ+QiMj1OiVFDT/VOHJc16/Mz7S0s1v/agt/g0nlm9S7nOv0saQU7N
1fevVsKbl+hzncNFkWwAvWjpY6Ncx7mqZGfNAzbnLaL0JgkXxAJM8kOZn9N1Kujl
0zO4NasDze/rurqOCXh7xUiYm8jmAMYZLAEOxczyMeHYBJzYHbJhfm2VHjSB5bVu
jgMP8IMLVXyv31DkmXihdvUZzPK/8sE1od/cu+0vJhY46QAcucpNviYFZDAJ5uGL
FfWnScpOuqrmq5bQU6l6QoTeu642Ldp2yA2rfnL4dfOV1lAW24aSd2aXR/fbhiFL
hQB9ISPI44LSlQpmeM5ALe6tc3uOFX/N3NlWnKFcT8T9CZEh5dOUpfmB9pJMyGfT
3lUcY/IJin9VsX7cBoGxVnKIp6Q5ubdw8lTeVxDhDmibMYi+e+nwXKQ36S55rCkU
5VXlmZZa1afTrXCul3Nt5Pmb6j2etCVkrw2a2uUy/HT8ViwdCgFb/N7CX+Y4gwDw
vnKMKmOOWKnOKJhkiUm4ahGT4Ugr39SBTVGpgn7KsHqamzeoyU04VTv6ShBjXrCh
Sf9ShzsB8aN10xEp5beb3fq6OJFEKObAcuZaHhsl8+iubeDDjRzvegEr9RTJ/k9H
C+YhMJWwhYYBdNgrbbeYJIkvpOoMuklqBYpnVfugMKSE7AL1vPhHJWOMbT/MTiIV
Y7KnqjedbeH+Y71ATUB0Z5OyuWZ2KWJx8egWahgbyWBues6sx5CFyppFRjlCYSAi
HR5i5t9+NzXwMhkPZTldJMlUYT/EMwb4fzB8g655B7/2CKHYRnkUu7XktTVWFYMj
DTvAYf2WLDe7sNR8afigvMZxwWYQj3C1dDo+PBjzy9+77o4k9z7K1d5W+qlQeV8I
/0DDtNg99hE/ef47G6l4f4eTsUKRt+CziH3i5hMqq86+EJ8GTX9jLCYuk56hP6PA
CG+l4Cq1QjughunGXos0Qnjulj3sDnN3YF85u1drFXyKKgC5QUOPW6DhPr80wbrn
hIx4lb9AfezjaGOWNk1txEHMh+FYdhkMz9QSKsFjLZlaui6X82+vixfCJg6Qf4V3
K7ULobzCZwSUb3dgx21rhS/x9dCZuyeJsW3fYbtUYQYA/bDoT932EOmPutLF7rvQ
6qjxOttEFoMO/RraykkxuP7sxiG77Vkx0AhFyQ5bpjhHzPa8ZvC0EdaFx/BQN9sw
Oole3m+n5lkG4o6xUm4lhjoCbyibGzJz6XTbslshDEtYowqX8PIn6SQvnHDByBzN
cxTFL5Nl1lXm1gXrtuNx6ALilm72ulY/QiMTTBolToW7KogjrhxbekXMUAU0ldmi
ktL310j389sjC34nxjWdnxMj57zpjbfcSDPYlKOVD2JuGB3I/OFWRQ+eG5hQF6vb
/5+572FND+1/ZZNegi8WCp30j1sQG4dBcn4vL/u82aqKfCUme0ja3D9EvpQ65hV2
1Kl8FXlQTfI6zxKJp+x/pqwvh5Kcda1XY7+rQtHbmwfdlyAZPO1+Yi/SsKdPs6R1
BKb4DiURrNyDvFVwof2uSH03kYRBXxaFBriNfSH0OWY02J79Jp/Y0dKF8E9EH81f
ZvszWfcUxDl082qJPXNOkq8uwnOWiemRh0UJVt2jmnuc09SuIJ63pWnWKm+8ylr8
qft2o0Aurq4pX3eZQzjALbjLpP+jcLy4GyYXy8lS8J+P30FPY9mF+27Ihfy/OifT
i7z645K3tUg8V2wEJTkLWPgGLcSmEeWelSYoD9X000Zlpmh6sRtzMkuyGbSADzIs
hsGB8vEfLgLCnqB01i6lrL+2EL+D1yb640JwjR38ZHdiOnlxEeL65xmHmC6QvPJ3
bTjD0ByOCWibBtQNHIlyUxnTdqN/U2nxds7m3e2Qw1CbDiwGShrwh6dfpDA+o92h
y1xoVGRMsQ2YJWg02tCQPyg4jk5QHmNmC/tKCF1okcH/xa8T1p3Ur0/wjih3nT72
aL6wyH5EZYbCMHBipo+u6Nm/HqzAF+8tfGVfIPRefvav0SWulqyA4W/pKT20azxf
VZ/t3TT11Y13TJQc4fu05ziFckRZ31nKDLd5DMGJXJeKLpO1ywvM3csKvoTXPJ2T
JoeKE5DiufQ+kd8JitakZ1w+j5qkLpS5eVaMJ4tJ+bxzkXhDZ+VkU39EKOEfHv9B
6tFhKrqrZtLeZjroDiEl7cYgUh+JkY64eA64EAXiL2GOykxeluD6ovQwImA8/u4a
ur6/LG9fBVgiMuZpYFHt9GNSvjP28wr9VuRLZrgd1okjdWcd2wje3LUrpiplTtZZ
4HbG5z651mYnUnXy9VHtgEWm68o5jWlR1EKZ0m+tmnwS23J5wxsZ39UdmjGrDGcs
e+BZTcophg0tL+iOHt29Yzo+OeFySQJxEHWfm+RDYWx5VXUHBhWDfEsq1/M04ZkY
GrF0NHIpw5hgdztoNYJBmUZOwgnILKgr5mOc0grOSI7rHAIZaXE104vzHqn00QRu
BiV/VSl8ou/PL/FXSQRZlnznwGLryO1wAnyGzW9ibu9BAyI/VgFM3PU6jNNq+vIk
nWt3EcnPBxVckEDYm4h7Mr3wEXGIagueDo02ittRyJGpHOa8qSJ1PBPiltrKaw0z
8imdoSkkPx5U/UL8c9nCk3C5EjezlaiMgs04Wp5nQ8kyhEZ7U+JikmilmRsi968E
pEum92Vi2fRbesiAZAKPxL2YIzqlhmOjSu9QJFWxKbD9iKwdQyqB/uKiwd4FGuV2
MalhD2gJ7F9pV09Xcfaqvmx5R614UYFON8hXXKkwI+Cr/4DLftvNhOkvsV32t6+G
vLZc3vKcfcf52qjP+EXtiF+LycMVmQQjcXA0Y9PNBICoiPS8yBju8VlNIuTJ/KMl
NbCo1Xne6np+iM8muyXUJ2OYt2QSDqJhCr2IO1SzK1dY7Z4LByU2zU8LfNFBvoSu
TNRGeYFfXpWPJkGTL8vy53Z98haBWvYUyglBtu+OzV7H5p4ahNEFcD799B7t04YT
8Br2rDGJNrRY0KQmD3jixhZWKFzt9l3AeJPjtL6wPGQeHMCOU7nbgIzraPh/SIH/
eoX0uCKCHklIir7HA5Vy7SjzA6U5g6XiE5onb43iQtr/D6lvjZzSnFOfYsd2P+um
kORl9nxAwmRgWsMu4GHlTulcCif/tXQubcAo8w4nroN1zNKvIHmn5l6zBOr18VZk
vSVW24iyMoPnV3MKhmDi5HUesdsMRApAgGUdSLt1MdHKJ76eQdfELLwEHH0vRPPO
w83vA66UsQWe4ddT4SVyerdeElyRZ2NoM6Rwwihjt4LXpdKL6Jny7iY8/XZA5Cbc
hcBX0Z9MhumCBbP4rmxnG7jcpvfa3gnbd6De3Af0fe5U0WTU2AvJnEZ8iyiIvfxX
N3gAdklpchXIQ/BsvCt1UI4sv7PFNyqAiImblwxsZYJczT/bRUxOLK6y8CdtkvxY
C/B7bmvf3t6lx0K1TOU34PP5ZVQ04pAVD8RkrUjj8M35BK598uum6OmtmGkPqKb3
V4W5k5lAnbq5YWWT5BquSPVov3/GvS+fWg3aFs1FisQjdjrw6nRvDNVOynTibSlY
ZSK06YHhMjfu6tSe0y8iV8hn41iEucMHpw2DHCCgAnyB1F93ndayhCWS+8AY1/u7
SdydRV2OtOVOixkA7CFausy/5vrS2UMjtzvR2G86LnJ3NAI7zc0Itk9YmbSOfFG2
Sjv8dst6qlScSBTBMiyJWcN/02eEgLjuiSssidXhYwwsiZdWkKevY/m6/hCMrv23
SzGgUZOSoOXbBP6MhbyJiT9fMO28zbwjpN+kX2HWKywu9KZ7llVmLSKL0AA1m7GX
dhCisffS5Lai8vM8/0Hko7rJ3UGEocjj4KztlV2wRylNnl9Je5EukV2PR49pHsxO
FN/q8X8NWjKjUa6jvOXWrvQCwqeGoYwe8hNV8nGt9lWmu83WSBHC2ESAwoU8EsEC
/0PfRIyAGYuRroLwowIXT9MQAiAvr7xVJJUqkIBDvmimH5brLeHYbUhGg8SUYs6I
sLS/EMC/mPy8pCPeInEy3RAgN71TkTFTh/jUp4xNtd3k9sfC+q6n/xoStt0axBEk
c5fPeYu/jtji3ASO1OnnCLC2ckxCk4nburJqAonEKN4uYWQCwcDTYe2eWVL27yeZ
43B6ZqIOpu3vTAOXSYsEtHoB9kE4tDkykPyr62yYmSD9yF1oOSOVHpbIqBTEuAUP
cvhKA47A3JUyiqJpqEJabujgdcRJhBXF9WuL7aNGYWeTOVxbCYpuO9v9xEPrCYXB
y0vRh57Yhl1YRW7XjZgc2thq3TxFSWLa3ws6lbbKEIajBz0Ho1vYzA+WY2TxuiUL
MKW2/0dkf1w8N2Mdf1x0H7Xft+fKv/S4HSIdul8K/C1BJIxz9r1gftYeunKIfgD5
uEISF5pfKJ0gh9d8pYMkaeY3j7Tl5pJuyoBx768vpnUUDq+9e/fyP+o8eGINZc5P
b42LiAoYpLKzBv1xKgBmXPgw+eMmOLm9GHCz79J+2Wjd4XCYZ2gEzQJEVvCt1wGx
hxz0vZhSYwkUGGY4W1p+wsd/iXAAWvbiQeEVvcG5SiBGNGxoDBVqlpL8tuh7TeCh
6FbpSh59W3HlIUGqB7+eFMslE9q1GxQx7P95UAKNyZadMPoerYahFNv3tZcoQVp0
XFw9q9/7/SttxOrBabtglskGFftx8Cd8R6PQgk0eAYxhX5mQY44Emq7sQ5VD87i8
e7PDvHKwDPB/NvEORSbIzJy6+T5t6IfspYWYEuEOpqgkgv8saTywQYG+J0AIUu9D
umknifejuLel/azAikfa4MlmFGMaoc+ZObbh88uyKVqrGkM6FvvWNvgjDeN8TNrN
S9v4r8B/smZPwp+hyCDM5fixfiYae923/vhq++O0hJLZzOQSynJU3wXTiH8kkygh
ig0VXgCNKFA+5NQLmDuBOaUmcVqMd/RFnQApUAZ+lJc+DyUSbwULJLrKrcbBpRcQ
cjBRsMWUihvyem3G0HBg9w8j7ldTnJhHS1z6NcnLL6+2gSQn3XIktzz2wewQohxD
u3jfNFxNTXy7F7Jp/vLZLfuG/Led1QSWWs8oEwsgGktdVSBS7vqHXv2zFtIpd2kx
MaYt+VOMlDt4F0MzpKol1HQ2AQETXI2PiSs9HIclmfCdp7sF0o4SJAATsvGuyMnC
+bThGWrtvdMwhJZT3mBDfgyMuVsk/RdkF8OLXvo7AHUgoiB6AA9dmQtOaVHbhiY8
+Dw0zLR4JnGhJfGhkUF2QkQFj1X5VGvKZmhPeRBLMOPGHEbSuMzjSiyTAn+E0m4G
oiCMwjiurlFneuhzwfC2+Nr6BPpS9jnesNjClS6jw5BT6Vg2hE8n0CRJTz4lIs+6
s635SbuiEotg7mgXQibIF1G5yGRFSR2QZ1K5MZy4HxytdSyO1QiHKOMqxuWZRbGa
ExdBwA+NFjq+ZWl9vDNgNuWl44xZVRv6m0HBwIJ/sTuo7/Ud9iwxyy8K9vKf/URz
MywnmlOEts9jc//tXmEV5uJAjDQPmBZjmWb87U+/tUa4QY/fn8LwzlleZZ4zzF85
C0t3WYF8nl72MX8DAubo3da+a5l3bp5UyDp2uLSxkQZPe/a0hJLIXw+q71Pmzdac
HodNs188HCe5/QEmPfsHeNXCsLA9bxma3qA8oBLx0cIk6JqDktQFLPntLeyZSAlx
nUvOVJqxxUUkTc1rsfhgQulhIf48YI1Cf2ssmzmRnGvAIwRdzaxmDagtJPejHbo6
a8Fn73RsXuVzrHRJ17ZH/EW97gBGtGE2cXIdO0wF+Sz1o0aj+G33ysRzSwkt3qCr
d3/caAuxDaWUv9YkwJjeKX+8+gVeNxCjfhPaewm5H3FEdqp07qkLp55F8G+baX8a
N+BciW3YHYORhMosaRgGVpa38ZU4lNaggKeX3+MtxMoE7c9LAQSFMB08lpprjLJB
xRaIgi7M9xbdM5T020PIv0oRxnpO/iWv1dNSoMYS+8EW4lFl2X5qioB6Oe4t8Na/
+ZGc6St0DSO/tpZwxLp4+5e5ZsA245w7qz2tfy2Q+gH+rufF86I4l7Bs6D30uEkP
n2m+jyIoUL2BeaIsCAKLimAwNhtDoOu92FOfDb9k3I2kZ0QMjuSDnW8t7h5YXwkc
4K/0iDxn1gZbBYv6dvEaWxDrCwzfI6OUGxfxEBZXQ83DSlK/JcuXElE1I1kyI8Dl
lO4Ybqcz+Sav60sYEpEJbuADuPwxjJZvY/66DXdFgYkw5qpHjLh0bV3eXVA8nhKy
Akyc86j2UQaweTyUXamtaPZJQBm8R2uR+XQiPWz6+lJPdWlR8CjCLczu+sh3a6iF
hgLypr56rW1AqjG17eI7052X5JRc6Q4RjYePaZrBNs7978nmJDfe5z+7/VFWTfEw
ChU/MmTkflritIuol0GuXn5DSsIqB3OrBX4saWWd8AACB3n7WLL3XqKxpM+rD+Uo
gQWLC35PcvXxhxjPsXwMlgnMLthhTDEdDl/TRcRlQv3IKSJFPRLlVtAy5FEIM9Sn
/gRLioIW7wW02wMbV+ZRaz3XhfHsFqZqdBIXuwQANjdUBeK7omPpZE44jpY9abmh
ZLqdPBHdqnfCHczY3yqM5Am+DLWfCnV+X1rPPwoQ3kuVLGcjrxFKAcAIfoxSaj+K
Xcb1BUYd2FF8S9KkNA/iRRsVcKOWn8t8u+ff3iAiBQr0Ezmqa40h49c1Mk2Xb7BJ
IxLeitvsFgrpcFJS4fYCi/4qCjugFkm+xnTt/tF+C3In5tCUTux/0aCcPgdrjuBz
BefuW899gNiUX39AJyT0Srb07gGhuEiT+KQB2QF0uEs+jVzsisCk4rEQLCX+k1VH
YHO6dTWpkSjg14h2oQPraZ1ApMEh21I1dGKfqmw9J5Th1O4x1SycOhgGOcAWDthf
KLBJDb/ZnD3N2JGXcpoQOMpxAZVKS1rTPR+gtGeS9o0yKgsx8r1xmAXo+ExzJznC
IDkjOZUvXhwPD2P6vvHIML9oEu9qsJIy0benEnwFPrO1RF9Y7MqK3gjc2q12xiFi
f1Mxwwnf9wyXFqD6XWY7+nsEvFtc4JVGFadOOxRnntZhpBy3n3vi8JbOlnP696I/
yUnIwP8OYCP+/YL0lDzNLW+cN3mHAHlr1mik/mRmMHqKCstIBG2L7xwxAd29a6Hu
y+LkMAlp9o+6LEC+WuCsRf0AJgs/OggprD261whL4oO/2KaMveVVVafmVfBR2UYi
sf2qiOvZh8LNNns7qkyVwEHPVkX1615GE+h6dKvS7/kGfl8E6W3OeGUJddttadKX
p0eFeb4Rt6oks/cQLzSSnLUNOAnLzbyQLHOJVcUSOa28KiLkInDhgG1idmHI0xxo
7LTAS/hyLoi4sHu99VQOcXvnzE0qdB0M+m699z9HbZ0Tg/5exbRQ9FTj4yrmkbB3
lFtIgeKy02gJrTOn6UEVk8WMEle8XZqkFYor8sP8scP6OltxCpzRyk2nm928nN76
0T1v/EJlEuU7JfgETggPouEW8v17mH7lSVKLLWK1kdUoI8Z4/Yxwvvtr0+s9Gdhi
oxVvmE3n1MFAME6Q0iFo7xAM+4FDKpFQOOYTDjPObxlH+GAgkELxcKAaRncofHMU
c18RzXx/rUTC3MtWCeJ8NPlofU6Rv/hiUOD2PkAuI4G5WL36NN2kTu+R/7bUWpoE
pR5Xv3T34LFakzle2YLmo6q3bTD2TdB639poZvWlEjYvUlyFIeSeMNJJcLmjwB6C
SyAYWFgvUp7Ai+pyL5X9sHvU4WQnEMtiiibIuEcHR8DYMcfzs0OaN0u/pxJf7zDU
zFD1k/PcvW6U1kFMbdNdmCPAcVdsU1JLqN70tM/3npK1nZnUSqsU1Uu25PFOUkPI
txVXhvH/maeT91DP/oBXfSLcDHFsvv9UBQn1OllNkeYwS54Q4IEsRtZAQluCkGkt
43Cai87W81OboSMbmXA5ZqARUuhlqM5awYKWqKc76wF9/OScgep9h6feMjxd8T/n
GepObLrCtMj53EFwYXLljnybLJ+e9WS0DZ/gjttPz19uxQMnjvHdNVA2+SLd72hn
7v5h0r9CqM6eJJg++pmN5oXCUfHBgi1WxQnP2q1S9yGeOts53A10cAMEihJ4lm1Y
MP1Nwe8pskDZRxqWUdrzHjLvuShHtlAbBF3M+ZBpDxnnQEGSLTu5d5HB5giNit50
xPpj2kxApghgjRh8cgSWMwJknjMrNJTk3PBE25eZwX/qIn7+S7oOWIyPI5V16cwQ
pcWKSet7eZs9+VcHd5glFbdoE9Rm6T5R5n9lF24BtQdaAUVngdz7oyW8D1SH16fk
QqGE7cYL1I6R41O7bUX/SN30g0r82h29iIczs2okh6O1RFGvGILa5gXZoZMsRyoO
yy6syTQSiBRp5lZ09u0JFyMt3zptaycUYmx/HhoGbiPUsH1WJYJ2yl289JG4A1jQ
IogcEA1vwU+IjQcfTXg9rfJ6NK5n2uD08DhspkDUBfe6mrs2ssuL0aEOevx9iuHA
2KBSoweuZDE8qdBxQdfYxmP7AXqwSVBsV3Q9abaXP5kH8IOue80c5DXGyMlJ9X0K
HRFJI21o5qLX4rH7psgbBpgi15qsiWD4wFExwrWLgnckpfWOMX5ux/eI2RkTEANI
KNzqAQzkkN8ed9iK4fUbEd3QHlvkd0+9L69D0rDWAQIWwdd9VKxWS6murClZZFgV
OwvQ9ucEzes5PmFg501ReK1qPEZmDKNAccylAb3vbcTH/ualPJp7NMCW6oOx02Kj
nhlU+pKtFSvB3deAmeKisaYmoIi2bLrHLyYM0p+MvLR5Zn/q+ZBUPs1boCQVkX90
SSjUYVeLKykiTOFPqEmG4fbxJ2xGdHj8vjoc0gyZ217v+xO939RMsRMOvU+OfpO2
OnT5MTp/WVEjqxJ6Ye+OSqeyGE8Rl87VWk1PP1i8qsDxKtlvbGehOGh09YaDaQAy
6p0fml7uEV1KGMKFy0DHl11wneOCon1+gJq0d0oQpmBXhz3EtosHPEy/f3XXhHNQ
MAfvRWYmgdMS0Hz6XRlqB0GTTw5csqmkYfcebP2anpu0Nozmz1E2HMhvZjaTtgcb
hz6qbj5L5fAR0muH2EF7pL8mTsD5LNistBWm66Fq/aZrIkcq32qCID8Z4WACwAYO
wHsUVDCqmXXd4H+TV949qt8HIdUwF19AaYblBiXIWk/tcMsPKSUwV2+wRp4RyHjV
Ody/bYYVNszGj8UcucaAh9RnzGvo7Y1WfmQff7zSG55DuarLXaGf0/5ijpW0SOOi
qJpt19SfTIAnnYgovDPkswt4QfeXpT2kOt3SD6UcLaLZLet/3KIQj4ACBmddMEMm
1lNubqHDP2E+/AC5LN9lSYQkHFqgBa5KIGTSMJifksVZqgSn3KdDj96B0nSsuZE5
Lm9mapaDCq/mC1tHiFvLLqZWKkvu92j2RIT3wAsKEmIPQHxBpPw1hCrMIldKdB7v
a+IbtOoP1PkZvD/aePkNdRd3ZAqorSWDD3xBd9GvZYq86iFRHxzQDWwa/IkmSWxR
qMa7/r4eh8dYx8RxzTM+Q4pim8fWE2bC2SlVbdMjYpcQtOf/soy7WnhBpbh4zGtd
ldvjm4E99a18F9RJuxuItBfRY/pha4jQ71MDG22QiKthz3C3fWWKpqonfnDr17Pb
qwph6ERJjaztlNy/ZEHvr3eIZMXqb8Uw0GmmTA/v4KTjzWjX/xsDuN/MHSUyThU0
y81gNNTzrcdHO+AxCFUJ1/H7jMjs4SjgboKVE+YdMkSID+h+cpRg2EVd9GNF1V+m
M9E9qNDumxCUWudNdu12SJPX+PitMN0PpeOxHShkEtDBnSyA1z6R4j5n12t2h3m/
D9ggT1qESpVndLzCNi0554VqE4mdBnKqo3OiU8mFnGERPbSUaUFAQkHKVaSsrWGK
vgqJjY17b3kqN16dhCZ+3krO15ZMLLtjDlRIA6ffjgV4x5kqiOMjjyOGeBt+Mfiw
Q5o63e1kCV+Zrd5QzPSNTmy6tS0gkNKLTJFoVUuK8hcY+DUWjxdvXuZVJNjgzNfO
s1Thzq4ReuyLo+v22/uoHYOCYgnnezjCfX+rs32CTQE4ENtVXEujbGtIXpnDQJv7
q0g6c71eCSRglQH+xZU5JS3VJjuCaFHRDW6yaGkdLFRZbx2n97YBxmpK/Ldc2hjj
9qVfyXkilKEvT5/ugf8/biQZnhP/hBOFLOQb8qTI9HE6GZP9+bQ6xQj2ju8XmGEU
6Xp68ctvQFX0SbSpjEEOCYyM48HYGt5Sg77W8e0kNNmYnppG1I1W/Ji7G0xdtzFN
hFpl04XHlQKE+0vJpoactRzF7fw0l6aaS78aE9f2VjorvbCMQXqng04AlOzgxG0k
jkHifAiF5dEa6b7/Xr7UZyEBXMM+naObsyoTT84Qo6fSfAogFrYWVfAQPj0zzF/W
Ady0ylBHPuZxYywN4VzPUDarkwTTcCKgharZCWkaHm4O0A1NfI6n1YlxCoXlq0Jx
nXOszGuaiEXBpo2dXXNgHPBPRderUPxDEXgi3qxuvwzd7KTXlJrPKNKJM1P5adMv
oHpddgo1CuE14/ZW5qWxw7Da9uWXjLtZd68Q/is3eXZ9N0h9ABHEe6r7zzu6hVTX
EEmXmOgeFjlI1amyklCPliKo7v7qFHLGDZ7uUrJBq+XcwuA4YMKzjz+ymrTkqRAo
8Q56RM1fcyBtL6sNmgd/NRzaWmv9nndy5Wcq/ngA1HYQiX4XEGtR7UFHiKm7ZqWJ
dY++N9UDKjzqJyLCZ+O4ncUJwcuOuXV/DFb/Uwg+qHajxGo3A3OfMYGLyqzbu4y/
UA7lte0/vOtXo3o+XRmbg9bYZxp5WgghTJSO0N0ZBIFDeECC+qEM7SlXkfecsluI
xg82bErGjkGWX4eRbK3AJRMvIrGsHlSB+32G0eppW67E6cHULB11aYNkWBSN8bLL
tM2JtXcBAo+k5WlWN+UCTGYicJfQXx3uK33DXCEAfxDvqdujAgA4pcWFaS1eYeys
s+XK5CyVkkMGj3khIewi/wUFcNzvvJRRLIwWr/v9LeW79tUEQrKBFU64Qd4y9Shw
ETZNuRuQ0S7V+Bk5B69SULPy0BAgK0uD9XjjZAUAIoTBoVxTCyrOGLlnX4XdDiGK
5lUZQKELheaw6bxPQtvC1+N6fPjesf+r1MRUP8jVUl/hC7qeMqr0uePYiFuzc70G
3pvY87EnrKw5+9K4yldWkM5Fem0IwKEvhV81dLoZ+OSuMlexaeMCMwi1DUR/nu6H
JEd9dVH35NQkFUUv2VkONAh4hlRcBQbyv0KynitiBq9G8qtuid9mANoZ/PVdMmHp
fJQ+hJ3EDHixIASc9ZXntVsCfvC5mPIcnSoLbgR68P0y6X7wWT3BipbGUPeVTdp0
BsStg7r+cwxGL6gXNittFLVY7XoWIcaZebTm37C0qW9/kWzo+bIcG5XPeJ0w8yHc
RrPUwXIFCBk4Mb3Hsxd6lCOSur6HSwzTxwV4UrCSk5SPpQitJdjh1kHi4W7ZOJdX
P61TmbALifjS1wxKpZXRb6HG/KMEl13tv72xG0JDhVBp0vNhTE+L5N5GFLpG82k0
4URtpC/5J0ONzg5gozNgL8X3cENynYzNlQTRqkG5Bl4GTel7Dgtq10UnwovMUBWk
F9jEpcSjGEPNpiU01t0cMTFJdO/b1BycEFSmzmIiHytv8+oPQRYlrE9XCcUTsW7z
a5+f9hsMdGV3WZawsTKhcuDQk37ACylD9CAc7Wwpz9ntibB1HnZYPtBZOFVcklgO
zgJvv/bM/Uge2hbZz4cTt45R1bug4ewj5t5SvH3ME/LuO3zxBHVw4iC211CQoaPI
8Pma32MW3wWvBuLEPpn5q/OwiETCxxJrpK0P7hcKEiaX15O2pO4QDazyo6JcyA1j
alRXuBir+XyTBZcvAESfGXgKSWPk+jcQ6Br5OrONwgT5oO7s+8P3eHaI784lU/mR
TLOj1RHMvYtKJovE/PGsttj2HubWpQWOFlMd1N27XFcYTb9rE2fqx/qb04Lc7nnO
Iy+SNK+2+kwgRpoI1peMXtrOSsAc6rlLOBtkBAggrR3kjY1vpNwce1B6XdO//r2H
Dm6LGX+4jbYWU2XGDWt8j2qcLXhXFLx8HLm+W+2aJqr6iIXdRGltCKIux+e1Klhn
VISekE8TGSfShszwmXaUR0EUMrC0XQsDHU0utmH7/waT1oZBv3QZ6hkkXOTTIFoz
Xhizvp18PRiGlB4ebjGPEziGLyzM4g4vmPUyTtIIjKEoHT3ur+XaNMlofRIyUbuM
tJfFgYxdFjvEDl/iaQOMOjNSB9232Q58C7vQq7LqX7giCNDOZB4nFoXbnPSWdZnq
ZGZNK1eW+Bg3TKCScCD1+7D3NPXawzv7t783tF3gN2kOLPFe+ANSdoQjkWx3i2vk
325e/PXLfM9sUQ17nh7oM+tJ7WL9AkK65d8H7gPSQiZHYTZVv3Am98PeUPtVvmKa
HVBiv8f6vliNvTRhXJOmNWbVD5258FMqzxgLEphgpvtHn6xlCEG0EhZIHwYOHiPs
He+qDDYGJgDENyzuoHLdyNfoFeWSUM2KzAlHxuEtlyN9xP9RI937YaRx+fXWzaqb
aTLwhIbQw5Ve/xpBrN0zBHhcVKEttVQOGRalr8aQFOmcKNp8K56/pHD1BUfLh41A
6LHJzWwRdspBQQ7NNgbzsUvyWlzWNLdTG5WKF+9pt09GgOkxl3NLvXTP6GKWITWY
6kGBkcuqUzyBcd5dinAttJ6mJili3oH5NsoCAAD2ApM53BQEL79qdc8zff6gDBwD
gzvIwLSPPfJ9UwTR/11lNrlzIZQViL+BFjBCe97w9zEEJqNpivhNYGiN5Zqn3HTD
Rm5PNg3cEB2evY5FdsBqbsd0g7uIYiryJg7oAUYT2QMkHhywkFZC7BuxjuAPxATp
92uLHKIklhH8t6u+4/X2dBb0EPS6L800+ZQlE82RnXDdkejkGP6lBqtKH3lvqmpf
AJPnWMxnPPF8vH6mPoGUU0RXao+Fm4qsFyWJdr8ceHBiAkZftH7a2Ciedl2Z2Cuj
irx6v5SDam7m34VT5gQNVmugFTw82CJwZDqIShnEidJv/lRtaXWc7ah+pHhR6d2K
0RmVLhXhInUqdT6/w2WsiDxYgA7DQc1/PpGVusofu3iHfPh+PBtYPngS6nogoKRS
UQINQkyBpXSUBiEcmmkVVHGQWpjEKj3jOZExVMWBGJrQQXd6G5QEJWBxN+ugQtM1
88SquN8Gl5/LiBy3OVgTeMvQCwjVhETePDOGlClB4lytFzZDE98rfMYPwHwy690v
iBh82BKIYScu3T7OlKI2xlK63zHkrPFnInAE+zgI+BO/aO0vFlB8mCiZxsIF9bTZ
MwdWAZla8r+vUMM0CmruO63fxOO6wveBJJNoYBYwd24+oHYoz8dQZNVkklfQ4B+j
MLfiCwefgXjzT9OrDpliem8mrr4ySnZGl3Is/E5xDEmWWbPYRyzOTebH1jVh5ZqY
zbEK83nDllGzggnZI6RXyecdmgnE3hewzmr0/u1gf8lrBjQ6+fCwwwS/+j/J7BJ8
E4mDvcGXBj6IcLXJrTeklIpzfB39i1SqhjJDctLm3ksT/l3oFbadxdpt9mWi+wB8
EUUJ2EziXTlD5N1aiUGLMaKbOiad52cO0mL6HBA/CKgdDK1Dj2xunhlQMVKZuK0l
AzVzPRa16j+9ulT2UL2IEx6uNAuCMnIaNEpwW9rHso87E6wveUjEuFZKgtOjjHh0
g/3Nbaio5UxQfsww8BzOHLipjpT3AEDlG2v+ipJ610Ay+ky3DeXy14BPzvzmpWUD
8I3bZEM5u2BzlQcq+U+FR//y1Ib3+d3W9lZYaBDXJpbdGWZxCkWKhf74UxYReQpF
YzhiXZkvdqI5/08/QJmJ7lMlMz3HWFnrWPOr0lcjic1LMGTi/ibkSTKnmWYl3cVH
MXlPLbvaiY5VoCOkmMlNcm/mJ6ulWIF6eiRsxGFxNyRRymwQwJAPEpTigR5TkO6n
V+deHVqaFRiWZxI/f75BYMNQHHKilhHSsLTlJZ6gMyag+ayPhvGptsFzpCsKsyAO
IjRV6cLo8+dVAqElY9u0rH059A8JG3Awl9OzqaDW6EJuuPtT3qitHPRkpUmSJG/f
VttAxeY79YGUOl90J/KWruR9pVLOFJOqD0/L7v8i3B0YP+nUtrq4QFeCXHj+ykFe
HkpPTGXjDYrIQuqMOepURJubEL0dfaJp+ZHfPAFAV7UP07SdTmvpk1Vqu+e/naxs
//GcxOHWEJDDU8vnngheLgZRkZsRrHZxRaAcZ/bhJVdkAf4gLIW5lcO/kqp8Pkxh
fJCvx8I2KylP+MQj0bOMoEvgCjQVYlns1cCAUWfx4nyDRero7kjx4M+wsdYE0Dxo
MkOHBRQ5zJ/ViWYDFsIvu03IWosSFOY0ss3BIjOaGp8/iyRNsb2RE7uIfFjirdYz
bplqsS4KRYNOOCq2zkTpKkL6QLmntyrpFWHiNZEraqlWrxqbPQDG5rit7oeUmdBZ
wUQu+CImlUWcgWYouof/72y0MeDVxQ9ihYlBJJyG+62p4EF0SgH7yYkkj5MxSK9H
7NUrDwaLVbgLeapVo+JrmC/lJGPiPvgVbxz2cPMT+EiPjnxF19LfdcWj28RDIOY5
5qB00EBhPeE4BGuACwUq+jKFkX/mWP//2DH3NU8bBi4Twlcd/LdLFJvecdIYcV5o
PcBwCfoOjgRvB4c4uy83siYzgYQkbzEZStM5YiqsIUefGa+xvHsMoxhZe6MYbMRK
8ULpbmb4jVQJ3WzPJs/LJBvJM9004dmpR0rjZ+oPvlOOvxKeovuXDBMRsHlotJfv
RZKLlU0Q5Wf2+bs7V5TcHRed6gipMc0ZcMwRHZ7BsgEcVVnSVht5iBgXCuSPHRrC
lcAv6OUaHkHaJ83diM5QeET71ScUlmALnIT+6UEMC8P6V8rnyErn+u9yZZkMCch/
zCu2GZ5bBJY5MmKPzPtK3BSzNloNpro0IIdgo+5pgHU7P4mywbZ8K3Ks2/iy//24
TWsACeqilqHnESmOKRdWI/0C8+s2a5Hxq6jSvNLAuh+Q8HyK96AJIApJDPpbPrXt
1bffSmlO11B5ZOPLOPZjLVlY4U6lySvKxKDlQc2sZU8c4lHNfrY3bC5/NrSjA8o2
j8TPaNXEeAL2KDV9HZR1Ya3Re3cpL9HpWYnpgMyE71O0exnZ41S7lzSZDj3n8KUW
kzJgUJkZeIj/zol1NLi9WJv1XvVj+plUolgrtVok5yO7Sz6HZ0pDvZUaaHczfmD2
sedNBREY1oQo+BeFBXM45mNj1opvbNMFZ0g+8Awxw/XsPyfo+qQYz3npeeDZ9l1b
o3jH6auit6g76WcriZ1mrGdC5brYtXKruwQjKrnqB19D/OAbXaKQQGBO9dYDP74x
kPiU04EkkG/PArgCFMDzckhOGQ+NCKfnkSMJs8rTYKR3K5JWF/5CFj8X4MBdUuNS
qAv0PjmV3NWJAG8RRNC0Dvlwy/xMsfY1fWkHpm7+a/tw9x9Es6ojRHOxYknS4317
vM4Nltsr5tncRh4cMu2NB+KOjUnnsGjkZ7JxFtQmLUTth0qmqS38Y8qAbxbYRR/v
RFapQnhQ12IXw6Nl4yHCZTQ+pd9mcT1isMfGMzf+bZem7+w3lH5Mr/4tNwHKZW+f
OTMVqfw+TChOsF5jhzQDzonPDHyZ8t3LumtiGDVLIRoZhzoK6YgkIWHjTOtyowmj
vVpU39JEcTntGSiqM7d41AWcl+ddgPEWJGQbClvRIpiS9348SRGko/10JRWWUEZr
7MONsd67Ph4t5DYuutyox2RlDp5iTIah36PVX2IzK6fXi18Yby7EKEZTI4UTRvbm
Mqf54RBoJmSFVKEynPsfk+zPg180lp7a2+CIqWLuA0cygkjhWGqLPSgg8e3zviuG
JzBhj6eh//nqk/6BMDOmfUeQte07H7UrcNhb6uzmOECargS2/OQ9Seyzwirg2ojj
8BbZ16OW/eKpVkpyAOR8HTo21D4D16iUq+GhlBE0UIYS1COcMGi8PHKIfpgDCtue
bMWUqehV3mpmcyLZoVse70r023xbAxgZdr6RzjD++C/KP2uEpdUWlh/G+JTtvzda
cX3tEyB/qYuXns13GE9nM66RHK5BKzGMpvvxqcf3XPhQ9RaKEgfMqcBV9Liq7nVK
qa1k52CrE5FFNYL2wYOQdK56dyDd7mM7LeEdTq/6DfeIIgckQsY6jlIgHilFnCrD
WxPpOa/YrXzn8vuuUK+iqOdovL9241Namj3Wg1RzygnvTndP91XxIexMwwW3iAm5
mQZidyL3SBclptrcOHacpugvQYiNbnpcgArBUOyBAk40+F+TwklOF0UQFhtlHD+9
L31dTlVMTE3QK79foMHUXOB6ZAU3lprq1+45MBaVz4iGA/frTPTNrRoFOAFfek0j
5uL4NCOoh3eqAsgKWVdeK+PKj1vCdppUfT/zJUhCYKnggJj41WnmyhzyciTge20d
6PseJUOr7ucn8RIJwS5cFGb4rD6tMtDyM0ltXZBIp2fPrh/Ca9G91cka0z/0TdT0
mrcbdVc8AKpxBV+4aLKN87sOZiDuS5igTP6gEwVBXqklbH6ntQ39uYJWgyS1ULlK
KdfQ67oB0YmpOlmuJyIJ3zSmM+5Ea9Mj3M+MQ4y4NoeZOvJwS7qko0YjsA8NWoq2
Dno4NGU+LiJU/PXBD6evnP99GximnRTjLbzdg6bmi/0+1Zply8kIOovNBVzFKmGX
elGxt3TlWH8fox07uCuJQYICmVHWSSqlwRYhRcRB4mbYLVr5PclhOZnVLe8cKCp5
ENUURI0U5CY3hxqHi75cf/J0KoP39j6aosB47RQyIk8/BxVSkwSjpmM8auzR9k7/
ecX89nFLoMHHByigIPDq2NGwIJiH8kzv8GoQnHRiCAbuQByvjIyp7AEbH1/mCY3Y
7JHxeMTN7CC7R2Sg+Dt8v8gi0NcxvfnEk6RRr5PBAZPFoXsNuQAJieVd1E0egND4
535WJt2TiK5y4WhfTF5a1xqBkq80K4mnz/WexBXrn/k/DrBzQtixbSeGPUuWJ8OB
h/aY7/M6IQu8seMPbQb/Sp3Ip304qhDo9fBIdPEYbFAtsVuqyBA0tAmN2jk7HN+D
L7mYA6y/5AQTTK1MwvqARn7Hule/IosdYkWNhDD4zWvvl2/2A8QkUvkDHXISu7um
THZKKXMlH1NlQYTgLeyTk9MHQtGAnakppINFoBExqBd1z9qvEkvI9ZomkJ1pUQXu
xcwxs5KntuGntENP0/YCEWX2wyyLvIiwCsdcpzu1kiQ88Es41Mk1NZWiCpHFgOEY
vDWysrOctsmS13YU4vtFGdxbnjIMNM91nJ9QioGueqd6jXRPgNgJ0yqfeAzJwXab
k7IPSqWh8d+qdHGqdLntYAodaiYAxfdZJ7XnDNfnT6Nfa7BO6QtxVmGrxxtHLtY1
l/ACwOr2Nunq2x8e9k1ulXF0bWU+FZByI3cetuzPi894zma5lSGOgTJIdd7nOVx4
eWU6FAvLQHRkZOZ0yjDIRnDP6Q14PABA3dBckrKMcL8UqZCnjgW7eewsrM05g+e5
0qIkuumSs4eX1FzvIJgd5ozqPYqy1tfUaxCiKU8ES0qug3z3O/v9DDqad5jSpFNq
Kns+LfTT7fLko7UMDXeuRNJpTf/hsUFiwpi8wg9+3SN64XKYJa4CHU9p7jTYaUfR
ADggG138ZLcy+ZXyqxu52+EXXbmzRigsW6CDL5g4hL1VA0PsgsuZ9tZZ03J/37IM
0FZd4X9qW6ee5RegRu09C8OjTQspMRDnpVSGmOYPX3yk+NLZUuiL+mB9O8FJy1Di
Belk/Avn4lfLS2YVwSuhAH4uR5Nq61ruklxiLbSu23MsfAZKtuoV5911f4R76xRe
VFkkE5P2i3z8ovS1bukZQ+nBjcMHF2IdBYvbs3YEm7ziXQl8emVxdlbM7L5oc4Nh
ie0dOzRFlPsNcGk2PhxxmWnPnNK4R6WTsFt/FqPf7NAu50W6+OKbl2wMlcE3YBJd
h3h+RRc78W8IKVOAiFyjuZvk48rivGq/qkj8RD0D3CcNHb4AkMaS+vjiU3wc/cI2
hrZ6YPhFoJbpcS1/g+0aeyHF4zShxfsbRPn4TdZdfjb2Tt01S/+w7dpt7XOogLAj
dZqzmzQXPpyk6re7vvoU1SwXkXGGaOxcpAfymvJfoghSpUNN6gNADLQzkH0CSXUr
EaLhpFMs/QSgSTrHZkiSFQgrqmgcmqqaDH8QEAN6oOIOvR//FA23tnZK3ElcuwT9
blK7kI1WxL38Nkxfjv/sODSJaye8sg6j3WlQef6Bjkkz1FpQTbBVHEPQXIO3KBZ5
9dSD8LKPPldFZc2G4UY7mrvK+1TmP8lV7eop8ZIDUDVpMfGj/Ff8arYIzjDLnrd5
+S+fzutQpGIelR68G7cz39dLC0Vf4Muty4Gh1X9I6CTbIvGq3dhcerIAukg44gE2
CzvcNy4dU3wosCySd4hz6Hor9o84n0JJNNat4Nb2KKquPluC+UYrf5v0RPRRGGqk
9j9t7Q3aaJ+urXwm4y/3TQREkF6tp5Ifu1f2CozCMPQd55qrjamgr8kFy+j5P702
w7/0/ACGVuxKFrrO1M0h1EM6x+S0BBJ+Jnrl1KDIqqmLs0P71zenTuU+Hq+VmwdU
RRjZq5Uyel3b3tXrsSYmgYUfSGPhDCmGeyuzPC9c8f0VL7wRSJ1Fff+V0ChDoppz
oie6prSAiOkE175ic0siv9uwPxQjFlPEOjHeJSha7UjanMFO7ObARI5KkDy/28jb
Y+cROyLbL07NhP0bIR6Odd1qG9hzG8TTWffdDSIU5FvNsP+3VYttvtDLcaMXh+Br
+DEkBsaP0MHSm8m0oSxM6QIXmRqBE7JRKrZqLCgp47Py63D20A8cwti5Vj7jGhiN
d8/rbDKwTPjhgUCWRa8AXfr63pAzktf5qUbYZidMic7Na6b6OlWo3fHTjts+hN05
s424p/auS+EkZf6ImAkA1YW81QUHwqGjjE3F4hXAFb6GeQjGglhFDm0UNefKwJsp
9/y3C6B5zuSPTt2G4Etqr1u1ZSPXUB2lPhKn9R2HMjfi7MxGASlrC6B8tOVExA9q
oXfaOd6nrwiVrvTXPw9xEEQnZbcYWUp2WSPtEArV1+hX67LE1irmi5dg5vDuycXz
Kk3ZmMvPqZsi33uL/h7h2UyRLZr+ZWgGbRsYZAEgRx3feGzd6k9M4VNwVrTl9Dx5
aMoq8rbCqn3KvSlD8M1U7XZYMiLBM4+UA2oYtl5wfMoUYij/A3wy5ibj4X6+ahtw
Oq2SbAS+bdDfWE+pvUwNbmaFWDyO2h2mX/KQMdiCd/88ZO2HI0Ih01tLIwR+8aLh
av8pm3sdgj7R7VtylaXZed/C0Xh2W8w9645wYuHbQ7SiOriFMKvvqlLb3YI+0M4F
8ly3IGPFqZzWoUXqu6cmTOBpgvThZrBQsSgc6MAmBv+FHrhOfo2SGXVhD8oBTfez
/j5Mjyk2rXI0C48uyEW4hS67ikjTHsdJr/scgzx0Ods99K6DWc2Xdpxve+BEGnMm
0H2McJ+8cChsP01EO48qWhF5UHWl02g3SUa4EGLyp+Dh0Z0he/xV64orFryCC12m
O3E2xP3c28SuBimHq3gQYSDUFB7/hxwt1i7O+45V+meZ969mUOgBCRxk5VxR+RdF
F2ywCQ7N63toyYOe/RClo8pq1R9ImqUDOvjc89AAo7hEDZ1xiJ8/cuLTu+LbS3e+
B38AaYZX9orBxIoeaa+snq6W5lPZhMOaijcPdkXneaamqi6FWN6d+SkT41giLz8K
kRe/2SBpF3lqgm4V9/oJqmYGGf8FNcQpTOh1RKeLfX6w1N38gBDVMRxs7126jDg+
z/fjZ1N3FxwrrryBRArwh7LEnkNB/LW2h6WwJ27eQf6XXzJHnV7pPGDNhpM5FIha
kDq3xMwKjTgOJELBXYrADRmNyhYDLWZf+OBSA1BH0fe9jBPtWWfn4fwOvI7GHjoo
dM/j8SSUIvFPDY6TBmjz9qsJEOmGKgpkdhroWur6nNJd5ezsQInzsrTewZHjR7UA
KZSHXY3+3zFk60xn+j86DYjqutYqbz6kTMW3Ai5CHFlz8FpgLAgoMqhoaIuB/XbN
r9x4mCIIxcPO6czDfRN4MrS//cJe4qkNP066FaU4/pMhDPYt0xj3CpBRV4GFuBZ9
pwREyTKxaoQDT4LymvCbUpAnnYWSOxLTPpCkS9ST6RFU6WldAaracHb47MzG1Z3g
8kqI1QlXhyUZ87hy98jqZbybBctS3hQFd/w5KktuhSK2RXJpPxcd7GLsYErdljY2
DFD10QIXltAJy8WGgc3n/q0OWw/C2uudaQzR1Indf8XBt57Mqkq+5g4XIJvCr3Wy
c64/l3J3xwCQV7IOmM8L4DyVY6lNdvTpzIc3ckcXT0J6MHuy0QRgtvHx2ks487WQ
JLhrMMFT0Eow0Nn23qw9m+t8OjWsToEUkogg8FVlpoeTcvtrMJD0DQiezIY2Ae+U
mbzocFhgM8IR/fHRlMDzzHfCQPVAHeDRvnlUaw4v/hhvT1F/s63yW8sUICp4NDS8
P/Dx7yganbzEsJer9zlUrK/ce09dPbrt0GDklwM+QGXxh9MZLAAUaDm24L+Q9ilF
ZpXVQX6u/B1X3CrqOnQU/7pHHNNiQApzWbMbC5or1areVSkLiEK42d+zPUjmMjjH
xS6qX+7eP2D9haL/4ese1OSDELIokCSBNONpnPKW4UfKhcCtfidC6TxNNdwiHIl9
84SlqTnxec0KwdKCSWlwf6ElbZ9ZZjWqyb/6CiJTfthDkdAYGBMXWApdebodI2Ek
/T7hUpPLiFfY352/C/M+BdKcDI3KWU/AoRYBCOfcVsnEI173RE6h6pmN4fsvEbIO
mf/o7nSi0GGiDa0akP+bMb2my5oozgK3YLLb1BZFYHkS0yBeI/iYju69khwWj62m
H91dEiD9pTzYvI8KwaQV5zAT0ul9LbIQE828rl00FZYUC4MsfW2KQJ5E9YzHxYs6
LYCF5yOVFajnWnwissSpvq8l7j4pffE30bMsFyvI1c3pQgXRDuoQ/DfoPkQqg0v7
iaD8um+noX4aC44ghklWuEY2kUGW9BUaKF7h1yniesB2+w/wmQHxZiBIuKkKJqKH
Q8Hw1xF6FY47ACynjogjWEoveoijHr0TyqjGNxqUOD+Do/P34aRzPe222/95ZHdN
srihh3gTtNTqsOkO+nc2PqBOSr8T//fk0A7qNuDfcxN0HPz2eHSoCtaKrMxNI+1Y
AP/dHWwMJnLY1aXsv4qNiwK4X1es7a+Hh9ixqBW+goFM0jv2WqmYb6oO4zXfnAm2
YeIePfFa2CNpYSyCUWehYrQN/ci/baooQ6yTHJSlNl5rhi4Kn1Haoxosof59uyIW
w0D/EpNd8E0mFhtkMk/FrDDYPTB8F/HFzJOvds4XFJh8n3RvNTAayAL6ujOsbCYD
xPz/MCHcSzggNcnjytMrZSSLcYp6cHpx+dU+dGdep6E/3kQpZEWe4YG7heThyaax
JeIBubNcsDfxXuZS72ZHADMiEi9Z+8tCT+hRZB1rSA9JutlkcbqAbevCeDKE38AQ
VxOfTPj3XwICwnddhl2wChXAT3BGeKt7oqF2UBBK8hdT+Rf5fdmCSnq+WDRi87mC
9UTWJ24t14RKwPbByeXBDYNg8oQpD20TMHlBVFyYr+My8ZN0LUB0lIjmAPscfewL
0ozcvUTwu9Iyg6iVb7ghgmWjmM/SPTM/LvxxQ5Pjuu5E5W9jBJq/BgF7+bVDqDBI
vhWxN30dgeoY2J8JPYhhFQSQkylGreVNTIohveCEMg7gISDG/LFjf90vKXZ3GxJp
FqoSsQX1uhBIrtfJbnkTxoX0AJqZE7zgt40+W18Ujb5pkJeot8FhBLZutfWS0T3k
w+l50MQLnJtcL8VBV25x2PkhPn5Q4fsYp3JjWzx8Dhq/q46BksElXpq1kdkQA/rM
2oV7dxd6qxOWcfihMMi29tqvgR2tbP725hBifFj8dRGdnjOeT2suEHJn2nwC93Ia
tFD/lk8CUYI7neGL8E2efSQTbRHdcOuMpxRkoORjRrklBdQsrpQ68ZIzPJZY4VPC
qbEbyzO+yfdhlYQBJZhyleztT016O6jm0BpuX/zUszZpSB3ED5GCe1bODnFPyAYZ
RJygVlmrbiFcvVFGng1FAMCePhDsVqrW7faXwVqggouqj90gAnWuZk0KTrPjUZYU
SXhAshww3y6AEoM6WRvk3uQu/MQkEke8rAbkUyZS+zkuKNZ/JhIBPseF7j0QNddJ
ohCnm3gWDRHLKwLId3KJOzXuyqy5fiaZcUqGZPuv7oherw+m75bUOYkNqN5AWZ4i
yuBpyJ+3quI33lHgmrzzKFvDmREl9ovR+Hyfv4dFn6E3MXji6yvThWPI9AJx4ftY
hJDsqybexGiJsjC65frWmfiv8dptmci9f/8tKmNWssXu4GeEHs020lB2HpBy/Eju
ZfYNu3wXpa/3+WGQq167c35GLQZqiJvNgZ85em65/Myoyzqc0c3XVGsL4BO1TZOP
suEnZHN5pLZARQ7qzy4ZK5EZH8FygkSa3ijWm6PvGuDz3PeM869I0AUpD1Xfu4Qj
EizerYbAnbKYQQ3s2wi87ouzjIWjG6gF2XMpxYm3laBgtae85PBjZccQLjcudpLx
0ubaKJSRz8qX+vNOi+NUIRI0q6eyF7UBnDgHVdUJPDHU5ROZLQ0zqrV46Egx45LP
eSYxQTCzi9sQ9c0beDBu1a5QBmomcdaC6lI2gy0txlISAGBZfHLwS/4wFNESxIF+
tzdjLZWQCKZ/342dieeDzbCQQZRzpimBIknsAZDdeUZAqoE9MnC5dD5SG89YHU4O
eSvKsoueL5dfezORlVu1kREdyEG8CIT4e8Y2TZZ20c7lSmQL8vcoCprrxOuipDf1
fw5EHeHp0LdFMQW8a3A8DO+JO6xidjeV6foBHvIWSxwBd5VptI14Tw6+KDx/abK2
43r8wyYGqZPJFPDESFRGybjFZvDrtImMBqMSGIOsBF5HtxTvj7Be7+Qv65ZqxwIc
/9+8ZExRvzQAri7bicTiIwh50Fu4+EhjumkKXcYBCG62MUOp+WRRTuLxRcBdIcLi
wXot4kMpRXG3ZOtwt8bGkKprsG+Nr+wUPktI4cVhk+xWEJGseb24YfQtUSWwHd/5
rOTMMIOS1f2xuH7SLpjGAZ0PeahoPMTyWrdfNvx3PUk3VvLw2rdrwHm4bjqfLDJW
yjfOt4846+wmQyMtVUm7ed6d9TQCPnkwQKdeck46qcacMUP929hBh1neGXj9bgNC
6bXnRYqcBnnlRzT3Sfd+Ic5ipIFOkz9H9XjXwJL5ge82FdzWtVPzKYzxVzrfMHHV
ZSHWJzMs64td3ikF981KiN1eQc1XtotXZfSufliMaTRLJqH/xgrpSDmpRip1thYp
NkYuSWmxSUkayD6SoFEQHZJLuE/iKdUDp4/khQIsTGpdIKmliCssDeh94FG5hzcE
OQqk/cGN1kW1KXrer30e4N8MX1+pUeOAUFL80STem57/Rug0ZAwJK7fXsy+YZqAF
KrIQZTWBBRYKooSdUM+owf3NKfj4Q60+qsgbJML/EYeQtdKWzaYgWIvmhqsA5AvU
kV9T3vCQXuSPoLe5kwaPzlAMiHNWR4NQ5ihEA2Ydy7yj0o9+ZJSARkh1/33ml1ZG
bSomZ+ScclpuDHSle3IPjO+blyi+/frTgNn+vHhyKB5xXK0yvBz4w8cNfS5x0f9O
jX79U7Z0lb1Q0ngGsaNoYpW39eapCmjF7WBRKBhlRGBoefMX+4fg3BJ+jIJpc6AU
n5q8GzoCrrY20JQf/qaeL+NTpWatw6ZLeSEW/0/5W+9pSGvh6ln+amifmoqqei+G
7EZE+tI77YJKfsPsfOYAlox9mpgRCXUleuffXF8yzhJelNJlQ6LGLIcZzK8Q2ccd
j05B5wcd9YslZriu4wojD2TBlpAsPXHzu6eECbVq8/brQRIUfTC5nwOA/2dCS5nz
mfO4vDONbRpD6rNZt+iq9f7xnivg7wHc7CCuHPknRhwrh8kXhRzGqFMLMHa+LLEC
ngjCKo3pk6QfMJs4Rd3fWHxTNl3g+Ej3LRLAJJw/quh3CURweuq/7Aywz+5zdNbw
nDjUoi/Z7znVEdl7W04zzqDcF1xhGuJl+nXgBLi855kbJ6TEZLoIn4RuuC/TRw+X
bYILSClj4SIGw5hFKxiWWw4pr0owJqiO8XSih9d8AfIWq5Fm9V8RYJEJo7ZrsJFq
Qr3PX50uNPkMpYrsJswmvl2tBRtBVpPAgLZvabTjmn5ASf7gXDFQE0NqoekzmHJx
htFFv2B3HJfUjOEtxAEMqJFiOriUd5E35THEquMJvPYeo4GJWf62rl4EIH3rICwv
l75kqqQ84lbj/HG0bVGRA63tYx6WXcygoeibs8+tY7Ocn7+zrgrgJHsLMPstIc4K
Eblc4TSr6ImHGUQzgyq1GpQRVGD+vtHazXvKvcr/5qpJ1dg0HWb8lGZGuORfg181
wA4MDori1mZ7MTkYfhMDZF17gvtYQTXabg+vD94F3msB0rqeRyYKG8hYSzUzP+2J
6SfSCd0vfkRtgJi4de1Vmzeh4s8GMfD5HNGuwxL62mS/XnxR7xHIEZ7M3o8AzwBR
7Aig8Ebr4e2V11pW7F+fhUwuGtAIEG4nSwiHQJ5lG037PihSjRR3xCTKcPsoyTaE
SVl8G0ubp/JZVwzgK7YHJuu57NDCp/kl9e5ZsZoypXTuUeMtYVRlmkXy10YdJjJ6
YovQTDgZ4QmKz8dL+8nvbDW0rTnJS+JY/enZ29oqEmjV20Fz+4A+YlDIm6oMC353
xnbMytbFXxe/zZSWNkMygUGOIlIfZaha7oWAf/9F0ReJs5der94R1UsObgoC7KYV
RlaOe/T3uVaBjZhEgdHcHg9vWVp90Dx8H4KYhbgY06umqs5rh6hBXxbVWsopyvIS
ZdCIBlxeADrmXxlpQgcAWYpDS0pmX9Dtol/IjnZf/ED47GXpgfX8DKsZFZ9ShFc5
p4coQhJ8KCe77of6PqrjC0vApLOBpmcczdkYD+0U/NiwvzD+xaHvOlLDFJBjnlp7
bxWIgpYMRXvmliaGs3QJIzv8Xs04kSn4olKaZnbmv/OIE8jQ0odMX03BlrpaFvzq
Ds+rCEKFgmkL3NHrg1pybUqdZ3iZadId2RDDvtymBpa7d4cZTHADJ/0UqG7FC4hk
utxePQCH1WxJ84uBRT5mydfhob+TvWO93akR4E8bWfDgEgXyOwpaMRMi+EUBWVjr
rpYVTdxQchGflhnxe9pQB/YvmkA03q1msAJkSXk6SqBwoapGhZRRrz4zHDUD9D1e
Ec+sVAZYUmK4HdxJAJEHFQEswNW1DZVXAPIigW1QrXEGvBbergYD9qF52wr7AlgE
aXxGu1tMot6URgeDISQy+ejTsOlRRPa01xgJTTvecR1bVRBRSn/AwU+9Y1BH9ujQ
jJ0FLNMZygEMj7tKqNaxvaDCd/osfTBGx/KuimUB+A4Mo0s8NrQqJLVBOA/yOr+V
QsfJnRwdzYqjqEHrDIUSHF9hR4J/W+8jCFWjq5R2FwgFGys8iJOk0gCavGwr0/2V
VvPiTr18pgLz3pyXEzw7jFLAA9hVeboYOATBmfnlClAwsatyevFY6mN9vuSu/QL1
H/Ia8ANk86UDz607F9ZXfMFipXBmZzAzfQiuhyrfZV64Z9AuK3dC0q1VGgZTXLxC
H5NEbIlPjeQGdktLHU3AXIIdWhi0xg2aidCeeadVALrg+YmcdHOaJ61HW4cPzh6Y
k6QkkXukxeLklOSOPLBz8nfq3yYBEGydOIZYYxTnaNKq0exwlg+WJATSLkw1BSbp
V0LxIZFYqwZQd0cqGCqE6QrSQgc7JL7I7zy7wdTBDMcINN4d1rqjYm00nXZMxyac
IBg2Ou0ePS5okO8eiZduKgN9BZerRGPUiDy9qz4IKNVhbNlOjuDIbJ3qds1ju96i
/FwxFGEhbHcsTbzDZBNIvQ5Ej/cLOvSfZLPR3R3Zq6b3rnwSdxmVwwnlEMwmbigD
3bG0uw0RqzGjq3fKzXtPozbIaOTNfDJM9iCCy/I5iXiqrORoUDT00IUU4qxPTXSG
BTUHpEvvi7g5q9vFyRtQdYcXg3rBRD4ap30N+rkLq8DK099ia3EsKUtoTAacUtFP
82qgECfV7I0hvQPeM2lNQ6ItDEku9NCvZ4T4i4Q6Qnv/LMUVDn3yeFTqt5kWC/q1
wh/5zOhFLJEf3pZEJ+86Gn1G20lY6lZtP49Br9deTLsd/C17RHx+wH4GUr+99023
LafFYqTORtOWUFVSGY6uH3mPdYI4DdCV1IDkbK4caHSCcrcNAWCONqo4O58h3tRc
aBRW59eQihDWfOzY80BV3jJuqCl7K0Gf8enKLBhoXGs2kuEba4Z33fV40rXEAlSU
sbxkQrI+neYYmJpbA5XgYL3+t1TPdnpYjK1AP9PEUKJA8FSs0LiTOptIhV8hL3x6
L7isKyWj+Ry/O/1DnCEchvm57eRWSh7NLRT8ofwzjulykj+FYZcqs845cF5jR/FJ
mR+qWUaUF63ns4qU/HiSMN3OpnWrKPTS7hrKGznEK4GVwdckzoLi0OmBAXeQFrMf
yhzcb+KgEbDpNwBjGeJuev/zdzCzC0skb209G2xehBXkhlrzdsSZREhioyfEXWIH
efqdacDYyJroGdBxi3SqRoSy5KvxHmAWogp1y+8SD7AWT8XkKV+Tl8jhY8RdPlAr
SUSVrrxbGl7FoR1Gk7QytHFJT9y0zOCHKD6f8I4Wn1DF4FPD3nsdLgz+gEJElB5l
e7da4uMkF3VR3RXg7F2zPn5XvVNl6R0bjlgxF1fYpdMhZTNz57e/ndLrvg9UFviF
q3Bi0jGTjrg0Wev95+Yr0snuDvRW9AeeQqOyTVAPoNpCbXt3weTkWTP6IQkabbbm
XpkvLNihjCB2VvDEE6adavp++jMud9UkkkYI8KH1nYHXTSPMOkTZPMuTpjDYKjIr
v+EJmUYjLmWaVJWRZQ97v5gg2TeQSJwPEYmt3zoBU5s8gSnjib23KFo+cBRig3h+
hiAbYsErIs7t3A4IsEA6P8OEDQmNtqI4RC2FuJT9FKD8vVbJ1VHH86l657NRGr4j
19bFDmeECLvkyM7bH22Dbmoo4OokCSeU5nzeMgr1Vo+wN41Q2XeCjqnc/nyBskEc
QxzquBMORjGl7JOW5PI1HszgLCG3CoxCpsr+F1DiJ49HYmRuzt3BGdioglRD0ug2
CVynm/qIKKJMavPLHxs/DHT6AVwX2OoSSGn2Rf8ob41wuE4IB0mqB0WeAKdyOKqL
r1nhQ1668LEuWYHD1/Kyo8s46RDANk0VJx0W6k7LxCGok8GIxHk5BQ8hdGybtjuT
TTJK02j8YvYuCHWeUJJXMC/7Ug0uqIXAiGcTQFf4NJp+rBg9fYOWy3XtKDcs773N
ZTtD1+qQwDTb4t0pCQV3op84lziPXmyMoUf1MDWvW7HOnRw3VJjRShoHkibyxx8N
dQLukarfVQqCZimWJXGQ+ncbfux6BeTaTL3DoPhDe/i36gbRYWKoFAEc9PnaBQ+B
iJ3LsmzxEB98g5Bs+KE0hDmDySYTifJbBRlq+ej6xpCABCmcEts4UCB18XmvhbxN
PMwccLTGAooJ84ifniPd0xiy9fXl1nHXefi9CQQNIv8Q0OosAmVYN9s2gZZApcr/
WV1lYpUi8cCRw4KGKPhs9ICeU4ic0zKi4FDNm4J4EgCYCl55sbM8fUyi/e9qgWuP
6BqeIs0iuhqwvmHqCxiSEw9KYVxl5TrCUmHMWJjECE0elFn4DzvetWdb9Aj65v5T
09ZSfT5hyVcpvL0UYH5QtWV1yuekWvH/q2zudrCoQry0+NF24NehiaNQtata3SWE
ZD0op41ohljR2Wy4X6PEBtDjnub0X8tRm2loPr3jSxsHJAj/QD3b39s6d1FWQn/P
YL70iAPMgZ17oc4/r7sGgA+Uq6SL4bxJR3UuPFZOfSFMUuQ3Pap0cWLl+JgMKVhw
fArbhNIX/czu8PWS2AxIw8jMiuy7B4eAvH21fxRPOPzWYTtP4R9QsNpxnyXPGFNb
taDX2bgpopC5bNTIR5zwwG0A3S2LYMtgL7JSVyn8DMVasiBZrAnj1IEFrVDWL6yg
gmNdsrFQWAs+XTmkQ88yqUTgRqzIN0LIDULvocXiltnkRNrCe95QfD7YiIm1BGtn
HaQ7mwLHOpGI67MlKK8PSSzWvZntqARfwjfhkrf8PmHK+JNHQ0Lo8P3CXC65IZvQ
go2rOjo8Zf55IFS4xfeDtihogXf0NBAQKGPuMU9OA4janlxkM+CP6JBTSOSW8Ayg
7cW72TzXEmzil2DYxEBaSEkWmub5xqdkh4ATtIy9LJ4s/aeK6wAIDHKpzs32pBdU
KY4ZSiOZa1r06Smbu/eMGro3BhsStzrzVc2u6frpuEBYv6lQ4icc7Nd8SHlDmSem
Y0wAYXUpx/viF0Up5OMJHgPdY6N9sMBxSx6FWDyF0m5bvqcGpIPR6U2/fgnjmg7p
/MTiOh2qkclohHyEuRLWY4cbbPnhBIGWnjaBLArEqeF1lWzXf9NaLaJcU9YcdVSV
+XyrvjWBMs1OvPLWzQuebLKO+BvHNuznKNK9jATIRApMUfop/FpRAHPNmO2xkByj
AK5+cj/2ELubzSsrrion+j8wfO9ZNo0IQ79DX7qSX1u6MsBOWAOECjDiQxD+kAma
vVqv7uSWS0Gp3V/EFgXZ+OJWKnYWrt3ggj6OPWNjl4U9pk9KHgdWftlR1El8Zqb8
RnOYnOQc0mYvS3pkNkDUi/qflGM+CF2HpMZviarM+Xu+dt/lSIMsfHHudFOlWqwP
2viAPyjLlWz6je8v2Eoe4vk9NBiTeW9iPiPQjW3Ji+5w2QAES3aI7lCNiOpkye+j
p5ICq3nfFNEEnKBQVpLIMe/4wCF19hV6Bb9s6z4xoSafqUTa5cfkwumuuGLPJ0LH
ySZmC8FlDWwK2RNX5NoglXnHL5TxhwdRG6xjkBCE0XwimmdyAi/J47lZ+Q4/D/8B
lCL/HLcpABaCDVbERQ6uCeYSXZ5l7nxcsMit3yyV8Ks1AYjToDx4RIqzWl5sY4mJ
1lMQgYi5wguPMOVRRp7KPP+LAdYQMHzzqb1qkY8NrREi+rnYzVRgK/EjGGj46vK8
BlU8XzrCGKygO48Ycf1quvLil4oT4B/0LEj5Y66gIhFypviEQ4tUbQEJdKfqg+GY
TAQBGX6aX0S6DzMCOV1rdUgrKScJfCNAUNibcSUf5bL8yv7ukuaBJZBsAQ2KQhV0
+SZipFctV5gUj4h0U8Lsq3ZuvZnVbmFRFhwxi+VNTnKco3mm/c3TXrZakABOq4m3
S8FN3oSfpL5RQ4NewFaxgdinFOEll1QFQGnnYYlCeb7y+a3uxK8tSraWGrc3kyZO
JkWdapp4iOnj2cEZZk19+yAXyQ0034a/qRYvM3CqW8g31GPVc+Lv4rxWfkFUjS9J
0ZNIsRAatXSxtcpi6V2xI03x3fzYE27idNQDO3JfhuQW8NW+mxTycoh5HJeiPXUP
dBUnAUfylr7ZkwUME8+7RhfS68fWPv/w3pvJnQCl7Tjx0BJM/GSktWytdBkRFeQs
E4AlzBOqQjUUJyM6tZmZRTEohd3mdT+NOWPxL3iIVGkVM7rkQXR1L3Boohv4pZdm
khHYeE/gFse1nT+nowVUl5r+AZPEi0Z39eO4iW0GsA8LI+K33wVuV9drVWNFMIIn
NKyRmWOy8Ui814KXc9b12sFwp83fKg23/XpL1Ko6IdYy0agYTuVKPFc6jejgtLCX
QHA1FcLZWDcN06x3pNlrcHhHYPjA0++lBM2DtAqa5pabEadGnw2/nbop64q3LVy/
zkZGVr12mnUDh7WfqqObxVea9slSlLg37yvJ2O67xkNe10ssn2YE0RLdo5Obj5+C
6UjNKLNxGUn7qFXGd829W5HCoszmwSB9vRksb38TonK4lmTgalifvpePm7w2t7M/
2O3K7bZnYTnPpJcMDQj/G6hwCpKAE2M+UGq9/YAqPzVzvyPGdp9Xld6GO2QizaVE
K9uhp8rI6io6Cs/jLk4irv0wTgXWvdE78hRVPrX90fVrr/tzST80xZH7AASBBwIG
v5xlIIGNTSHqqLX/0/3o/d7P9ysexYV7gckh4ujlnHWmEPFQmncy+FjsJbf8q8QZ
YAsEYaeVfmOiuVkvDZHMY8s0xyM0EjtkHnZ+NWKzKZiS4QbpMBd7HOeJznAjH1oj
Dd7co/miwrkrmFyBTm6w1dh74sUIRLpr6x9z/9Mec6KjSEhCh3Gw0jDD4S4PwlU5
KL7J2+0yQvc5idJ+Q0teoslPE5tTHI6/LzPcCInzFMrjZLwm9HL9Y1cSrutnVSwU
dl9kMLVCmLOuyyBdBhfuSKq07QXwdn4BNEq+NvYYh5vsj9/qarrqvpsgxDKQPDQX
6C7nuuJBCtKMkcaYA0UQBIsIYqR1Pm0+kuHogMVbvOftLncKXoe06+nI1EmT41mY
3GhLfjj2tzf1Meh/1Oo6GWV0hj52hkCUx9vO2JtsehLRiflngtOBDBPxCC3pBZ3d
gdC0q/MULVv3XHP9liQAsyFDFTr+BpnLFvlP60pYQupbBQpKj7uwxDOFrN8CSsHs
mScwsCEpPNUC9RvoL1EMW/29BLZTdRxWSQeXkokVRFGA/pJk9QItvpcUKdfgDZju
trfZ+Z/AK4IbHAvxi4sqjsiFZltiZVBfFvqhptW8jNebX4REJqQzqaciO7n2Hqqv
iotcjcZrg7IXqmZ8yF3IcJj151V6WPw7rmVZ6rblWEmxGb7ZYSbA1625635xhpfe
o+RyFqQOv+N2l2OtSr/vl3Mdtzjt59Z1wp5ZYATRuKpXYcO8GKloVYhz6bftmsBj
OLSbwfvWSLcM6f/8iXBd08NPWRPmYd9nEi1CQIzdO97k4wF6whp+pgEMPzgB4eX9
zkxCMB+LRh2+nFA6pkkoG813YeKKy29ZurZmuWCKnT3RQUu+rmg/bI32oBnE92HV
QQWkCCQ2Nw/PAQl48EY+nvn1qnoL9Xs9rIMLPMbmQZHdAVU2kBcGauVkCDcPbaRn
tk1MJ9V1W/eX3qZQfgFItjqQkZXH+BLupb1lY6dA+b3fqbHeQ8JnrWnbkV6+t3vC
rUGxbpJMSQZbl7NoMhLkRekaMmf3h7xp+gwMqxOn+Mxv9zp4oLiq1G7Q2ATx3jaa
yCjo1Le1QIc3fdSLBf/bwotWnaPrX1LqPHM3FDOE5LciRk4oLTE+ieEpr5frBu3P
did89dRfk9C55zG4I2RmxrX4rffe0kdi22orgaU1V2otjl5tYz1cyLQ4+0c8S7oh
KcbxmO3Al9qJqfKSUILot457JvI0M9ImnFyq/PJyvi3eQkOQjCR0wwSIks8oEkLg
RCRh72J4JEqb6yvZs4myH3MaoE1BmcwmNtTa5CKgMj5nZxP9e6RmUb4AH0NP7Efh
4Z1MVayAaV4l9h9gLD/6oAeKIjXWHUN2lS5R8LD8YkincmR4moRS4wo3k7URlQ1Z
jbjrM3PdFifId+Cm2c8NppBrxHZeNJScYTv68eC4vxa8o99I5c2wSeuw7L9pvzYl
nsYs4wgqQuT9SjdSnbEpvfIy0EYCp8eRiV5ajT2QNRATusDwu2H6flNzeBg74Y7r
+6LoU/09eZRlZUnGgVKPsWU5G2hN92WkiSO/wXO/kbGyhL7NskdelFx9KDTaVF+p
gor7QFxiP0eeQ87NeQ02hVHDEAOkJiIZG8ASAXqy7IJE+ZwwauF9p1h6F8brNhn3
WbvwJaqDMY0c6cUv5LsbbDMu1L3wpo6Ny7TYlQvjDPUDthlCkSHhO6TsJfDW2f+N
XLrdwv758MtsMatIV/aKqbOicjCaQPN7Lx6F8qzZDriElWC7P5PXxCh53hP1aVnP
Nd7wTy+jqAvHAcyW7mEw6zx6GnsMzP6xGTQopJ68gxhau3nGv1iafqTvashGgN7W
v4hq6V5PqNBKSYgI/keCvuUtwlqg8INWO1ZsqzPHcaaZLuJSLWI6VgrSeUILaU/9
xmwxOmj//W/2EVBomeO3JTUzwH/6buodgmRhy0sbsX1up/dpseScmfBYFOKhnf1G
9UEXT3lX/cRKmhpNP1KuL+gzLH9unfM3gwnt1NiGsoiK6VDj4BYHgWOcub3kcqDR
bWfAx1vyqUDZ6Wowmp8wH6gLKZFbsUR36RszIj2wSxrEGTTH5qpeWlBG4oaZAXcC
9ERGkQ8fl56wWWYyCBioxKWQQfdoDj6p2zOacBFD3xvICSnwGwYzGAaIbJiMLzbF
o0qJa5hwiDg6PYAU3rteDddMUTsZD0hQ0SRzxW2Ibjld9lCHM1q7x6zbXO5JY9ss
v0EUQYBoVCTwQCRNQGax5UkrEC8W3qcCgdlJhEpBflkZtD8AGPRJKUZl2/9Q6smC
dhR4Ldjs53qOcNkQaKC/HCXFuOo26sJZKnj6wzSmwafUZznolJopUjmHXYogtGgn
YIeJh23RyxONk8BvwOiYikoFMtSXSGeAiNNG6Hc30EUmmqLLyh1PvTFMvtChc0j5
CFA9Y8OFsgpQ03Zv06ZnTMIrjlZZu6uOLCUbUUlEPzmvsxcsMgN7WouJO8qE+qHe
EadyyvrZ06kyeNqW9LbQ8yzUA0uLX0cdSeQN0efbzB2aX3uCXBpA4UqbMxlkcuPa
rKNVuqXKY7NmYqJ12XgsMkSP4vbMGSrYAinA7wBtYbCKXZzZxR1rR0MZaslO39v1
yfp5WfeEK61ZQSqrcNamatV2EXcJ1DQKxyptTDb1+AzJ5KK8vYwgwTy3Ik8Fk7Db
ccY0u0VRm26qLMfLos4T+HB1diH7t9T09Sbj3x3P8VzFUwtGxmSclCHUy1vL9QjQ
XOs8/P1Tm7wGJHpMP3UOkpdR6FDcTW7geOUDg8VyvbBusKo5IyLozo67Bolkc4gv
Yx7aTjhaP4JkjrYKGkKk3RNDsIBWhyZgZhmW6vGYGfF4tk11XNYEm/PgrG8yx6XE
6/Qna+VJQW5zhA2pWa5znDEkeFZb17PwEYgcvBJWt00QFb6t/nnXoKj/LrEXAOVn
CWnP0SJ1u8VXV3j73waIS3S4FTUjWAS2vkFovtHihzFZajTmcyrnvoAaYFFxDn6G
z9FY0Go6CR/9yJNUugKIwk/2dz2P0TiFII7Hq5W02oBfp14/jirfMjTO6urhA+Bt
ryGCdt/dhaIsx7we3qbeFmufUHKYZW+p4Tkqs2dwTsdIqfFZsnsOAtYFX+sOjmMn
/ImjYxk6YJ7vq5Nc+7QKwrKBNas/XWle8iRO22WUZHP12qXm0I8pvEr3PJMpkrfC
IIO5i2/HrwUBbHadhhOm8bYkNlT5nnbg6yHz9HzGztvVXpzCU+Edcc9CxiQQxNvD
8PlEJa1+6nJ4kScqU6hOWbVgav36Gmjc/qM4cdeBv9w11qO+hK9ABzYgdvdOYzHu
Rz3UeD0HtMZPUGiZvFgl8uLuuSqWDqHlQDs6/9qGkfQwDaeoIEDkwpL05UqIBzrs
RDxlSjMildcKRuhnaDpLSxdbFCJEgPVHPDMSgPk2U1B5va2FWL+x/aeivVwcIiyr
BNO5zv/F/eYkKnllgO2+7hniran8Ibd3GL79yDHjOwtfmdZ25UW7qZaRttNOE5/0
SiEbGrdVDK7HgwE15d3djNv5kFFuCNEDXxAC9advxw4D/AZ8MbUwdx8mMfWYL7sc
wN06AhfGKJCHcU5JIiZK5S20j1c5VNeUPHTXC3rA15r0jio2i+jEqFGqKN4NtlVP
xkzCC8+hMN2b7JFE7CMv7hj6YLy2km85NmjCf4kRZQqYTYkBnBsIMM85DOCkgFG6
GLiZhXx71p4zjytCXSSguc2gWEotqie+EvFhVKEEjB1FbUbj8MA1pHM3dpYnbnmo
7/UzidHR9Ksly+gWKsH0hfp8lPsyunTDo+I5oN8loRuJo4b316iwxbi2ZA6wtQDR
oX0rLeblzhQyjBIMPv0i8EZ4V1dbDBNANlOUNwPFlzbGDqmFgBtwkCiUwMwtjV41
lsfu4c/kpT4XME6b/tCojG89wYB473aRDlk/wxfowMUCTYJ76gB7EGpjBfqd7I36
wDc9sNXap/satp8Yf7/1IXtFemob/P0NH+Q/K/6L1TjslvdMR8RNUmGPkgrbHt86
fAsnpjTIK4lInqtznPaZ8cf6AF1Send6IlK5IeLJTEiXg6gwqV2Dsf4dtcE+HHeA
AbONfYDOfenJmdY4fssvhDmJbjbxBUJjOCzOBZfJjYMg3r7msPuycgfD0/m4m0Eq
y+Un8IbU3g9ek8rTm4ZdpycmiPkU2Iv44KFu0y+B7wfoJf2KnhUejCO0wtmUV5SF
C6fuy6cuBmSrMb3MUzsH+9HaiKAR0CsQO4kb9PjJDoEqK5t87lcMrRbUxMl9RRAJ
uNZMxMY/QzGzP2hCftZbdX9kOWCbPAajaOWdGhpzu/qIZdJuwC8Sdh6DgWTVW2Y/
EAUrr/zUYPrMDkQ7GXkTJkuYV/1wE39mrz9jNpO5uGr9AtmgpGAiTusK3hb+B+a/
MHwhQTj8jTYv6wWAMD8LI2/22IZSSL4IeNZXej/CtM7oSco7baM77AFBoomBopf/
bficBh0AqgS969WPIlRHPyHGGizLKBFVMCGiyQx303KkY+JsMv50KPCARYxw/YQU
b7PlC8KInsRk9JKg8kzN292mORSdxOIwvf6yECLgr6ai6XHSDcNNYIlmyT8Yrmiw
neqEb7ZfUNfzVC2M5ncH+ZkBc1oQBCe7WuG37kcMHO7dtz4VfN59YB5m0UWOoTD2
6vafJdj0eYrwdLCvKQtrJwV/vUQsN7ZJctK4Mf3D1J7oyvxWwj0fAg4vuwzQ1yxl
jESFBRdPvgjrHBM3LqRgn7Rl1cjy2HmfqDyB/75AixPZcpupPQs4x6UbYO1RC0SX
W90jAclc677x0jAqgjUmhT/BGLpDGpS0rvkHQ6gVszsmdd0wwxHbO+wyUQ3PPoxB
SSI93VT2oFyLYFNvAZMxy6fINNw8DuCV7VGhubkGwMOLFb2pNMSaJvhJPpjHycgK
4Kc5RzcC7xsKblYwrLoShckOGLdBA9Os0pwRnebzvlh5ENN7p+ZjKKXgTjw4/AYa
qanWh4vDBeZqKPoGiG+JZA8o+ye2ThvBR+ekcjty1XfXQhDVzCeuj7DEqvLP7+ih
S91dOFMRsrw+GFa8RfGe1GkL06ci/1jwKawB7YJwt7Nxu7FYbevjUSZ3RUfcd2Z4
iyQloB5GuCkbD+8ExTXyL24sLezkHMw0jPkc64UD0Ulapwz+I/4Wg5Yxy+X53PhE
uhceQaWMCxPxviGRwUJzKbO7+xiGJv8JNp9b7HyM+KjyTlOam2kqNWCl/xefw5eI
RXi5TvDybW1U9DrAlCw3ByMO1IDZ7lu5zqJWOPRhNKquzEQfUG0LCsemjNOVxj37
Rlrbmf2lqI9re+kg5s7f7l3LrWOSrysyGBjBbHd37fqVs/jotwtg8+cB1g+oc3Fq
6BUyUurk3E3K5OETfXISZQrLUNs/ZnnEUng2lJtH9Pzg6ElF70CLLjIERKt4uXjT
9bAuOkh9kL3K20Jd9yV3oxc7nPIyCvZwoTFbOfa8YRNouf39UEZ3Ay+F6PwRXh5M
h1oiWS/wMPdknesht5EYl7hY1UBH/VhAtyo0r9MWoElISsrAcad7izvurxE/Z1Yh
vAqnr2VVNFJmT/Rqf3B2UgXB60ffzywwAb2ncQuamPNHfsKo1A+QAXkPZxfMWtQF
rYNJsTpB53WbFc081d14Fj+kutIgXuuwc4Ciyq8dHVmZgcnC2CKjSEy74b/PcNW5
QfirKjNY3+xcO5nKVr/2ZOn4EFbULjD8kSFn+UMFyQzJ9XwzJSBpW/z0Z1zSDnl6
f8UXf4w8rMoCHR5sW/YKqfo+RGgTgMbfvIjWijMT7pBu9PCr+nn9jyDh03umPNGS
FhCLRD7bJWUmM7u8JcnSGbiHfkZ2kjlAm1MdJLtCe/zFfgDeC0E1pO+WLPJFqcyz
c3ZbZTny6EP3tIu++UHT8dwUr9I9qGH12RxH2BYBWvqP5j1TZEGk9eLipKdS25c8
ga4NuVfb5ds9UHZmDoefeViED0R97f0wFUadDuiovp2q2z9y+uZbg5LGISyAieo0
RA0WaNEuVhPiZ0OuWNr7cxucEMJNYSTuhF3MoqqVCFfihjryEDg1ONi4bqKIUb5W
wTSCyQvasgefL6a8sOQFC5lvWVgNwJjJuhJYIcDrqO9NshLlLsTEKPUEEdYqeFXG
aykpvfROSS11JoS2akFjynbya0gxRb0MolWuDdb/imMO0zk3CiNf+X3inOiA0H13
/SzHwKTrNo1E0U/cLyhdswwUriBo4YlcXWkqYhrvjddZ6+WcPcYUmB6V7pfYsZnE
/Xj4CSt2wLUUT09PehxUy23HeQyTP1M5QyQHcfmCrhdj250TSLgeh/kcD/JfmlIC
LJ+ah6Mk6Wk8EkER6GNXn3TqTX12CpJR+OMvrMTQYHWV5mvOCfXUxWu9knHIJwDd
LXYJHrHH2KbWCxAsCVRnikCFrb0RzFRV/yr2iEQcR3S6epCXaDxsIryIGqKxBRcv
FLRCcAeO+zEdlQe/r7kk+CymXmPNfOhlJg6/H1U71JO4Tx0G8+L1z+i8b/5hUnph
OIRhuSuOJeC4M+ca8pLz3MWsCA/YmOXTzNrf+adgEYHqOmiJ29MxP9IYD8dv9stC
Pecz2rHqPMVnSBSJkpjc+uLDjft7l4Y0RJSdRPfjDdMv7d6mV5dHARG9JxolngPq
dSWB2qsPO6pV7Z+F/N/Ooe8fDEokBxzF0RAQagZxvGcyo0jRUWxDmSsA9UfHPz6Y
j158YrNo8zY1AycxW5j//AWxXwNc+/atpuI3ebqWGIv6dKKVs9Cs6VHT8vSqDRTo
DC40yBJlCjBQuVkak5w/+1hZkN9v3lYDopaS9SL6Og7lvfRWW4cl0e7P+Y59eLAx
fvcVUFX+xJIE8WvXTCFy3h+9KZQobr1Zgz1UWEL0FiV+S8RxdT2qkrZCM66G1GCW
vRY8sE1KFXYpSwD5S0rdcgiMVwEECIpOMRg9AbH02VSXaqcbtxLv4kWUsC09fehe
/Y28Ms/GHefHZY9DlDJEhHRT8byaO8tzdK8SV8LzQWTmySie+zib4wRKMivcI9ik
RoEYYqOtai5hFw4R6VM3uNTRk+R3URJpES2tieV+Q/O9FstX9eCcLWKYoSZQh4P3
1oFywJKcx4TCFHrplDU5wxHQHP/t1xpG+5XjaEsrYT7IIEZSXYa6iVylIHQNFEu2
Nwy86VwEyhR3Cdic3yNC6enVUSniRRmtDTor3NRhOKTkSvtCBO3U62SQ2saw3Isr
B1K2IJPAElWMLKF8RYr+ky9zBiVa4J/e3EBtS0Nkwl4moVESGv0B9NwhmbE8Ifz3
6IlWlyYveudorUAfY9F9EidTXcdWNibhUZXnRNxIgDDWdYUlj92n8RKA1GLe11fA
djCtDVJ8OgUkHQneQx7aVpepbbvD4Rwcib4Tadz46s5suroZyetKhwOzyhhFAyp/
9Z4Vy8ekgJpUN+dtxX1rt7BGlpuKh+4o6EvgZ572rbE5Vz+lLauh89T3CqR/B96I
jcz3vuN1QKNIiFacseAA4AKQ76TWLFGukoMHK2Qa70/IRJ1rB5owx8PKhrKT6Goh
EVllm77Qn7FTnJooo0xrkDnmk3LjQhqYa32SO07oLNLs3L8zhnSHtHZGR+9OOI3B
tSKmCA8nfXp4RwqXdkw+R52+P5D+7lkU26hgdogLeye7CEwzlOiPTyS4UDHunQBW
0cDgmA4kNVim46NXucg/73q5kriGGLDMIUmI3FI9HDRVEMkXcAahmVIkNV4n5ety
JTCw2LEUz68DnZEvUVkpYrYUhgTQAHoMoEMr9LsBHnywrj6p9jf0J9UYS48/R5F8
RU8Qi7+FCvWKAboepCiE/HcyG9kAlY5f9m966OyO4zhr05i7p/qTefOSNfcS9zls
zoof2RJPbeIox9aZwLcs/2rVSs4bLnwW6J27/uBDJqLSMOkuA1jgJSmcUQabtzmO
`pragma protect end_protected
