-- test.vhd

-- Generated using ACDS version 21.1 842

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity test is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity test;

architecture rtl of test is
	component simple_soma is
		generic (
			THRESHOLD  : integer := 10;
			TIME_WIDTH : integer := 8
		);
		port (
			clk                        : in  std_logic                    := 'X';             -- clk
			rst                        : in  std_logic                    := 'X';             -- reset
			avalon_master_1_address    : out std_logic;                                       -- address
			avs_m_read_synapse         : out std_logic;                                       -- read
			avs_m_readdata_synapse     : in  std_logic_vector(7 downto 0) := (others => 'X'); -- readdata
			m_synapse_waitrequest      : in  std_logic                    := 'X';             -- waitrequest
			m_spike_address            : out std_logic;                                       -- address
			avs_m_write_spike          : out std_logic;                                       -- write
			avs_m_writedata_spike_time : out std_logic_vector(7 downto 0);                    -- writedata
			m_spike_waitrequest        : in  std_logic                    := 'X';             -- waitrequest
			avs_m_address              : out std_logic;                                       -- address
			avs_m_waitrequest          : in  std_logic                    := 'X';             -- waitrequest
			avs_m_read_time            : out std_logic;                                       -- read
			avs_m_readdata_time        : in  std_logic_vector(7 downto 0) := (others => 'X')  -- readdata
		);
	end component simple_soma;

	component simple_synapse is
		generic (
			THRESHOLD  : integer := 10;
			TIME_WIDTH : integer := 8
		);
		port (
			clk                        : in  std_logic                    := 'X';             -- clk
			rst                        : in  std_logic                    := 'X';             -- reset
			avs_s_read_synapse         : in  std_logic                    := 'X';             -- read
			avs_s_readdata_synapse     : out std_logic_vector(7 downto 0);                    -- readdata
			s_synapse_waitrequest      : out std_logic;                                       -- waitrequest
			avs_s_write_spike          : in  std_logic                    := 'X';             -- write
			avs_s_writedata_spike_time : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			s_spike_waitrequest        : out std_logic;                                       -- waitrequest
			avs_s_address              : in  std_logic_vector(7 downto 0) := (others => 'X'); -- address
			avs_s_waitrequest          : out std_logic;                                       -- waitrequest
			avs_s_read_time            : in  std_logic                    := 'X';             -- read
			avs_s_readdata_time        : out std_logic_vector(7 downto 0)                     -- readdata
		);
	end component simple_synapse;

	component test_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                        : in  std_logic                    := 'X';             -- clk
			simple_soma_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                    := 'X';             -- reset
			simple_soma_0_m_spike_address                        : in  std_logic_vector(0 downto 0) := (others => 'X'); -- address
			simple_soma_0_m_spike_waitrequest                    : out std_logic;                                       -- waitrequest
			simple_soma_0_m_spike_write                          : in  std_logic                    := 'X';             -- write
			simple_soma_0_m_spike_writedata                      : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			simple_synapse_0_s_spike_write                       : out std_logic;                                       -- write
			simple_synapse_0_s_spike_writedata                   : out std_logic_vector(7 downto 0);                    -- writedata
			simple_synapse_0_s_spike_waitrequest                 : in  std_logic                    := 'X'              -- waitrequest
		);
	end component test_mm_interconnect_0;

	component test_mm_interconnect_1 is
		port (
			clk_0_clk_clk                                        : in  std_logic                    := 'X';             -- clk
			simple_soma_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                    := 'X';             -- reset
			simple_soma_0_m_synapse_address                      : in  std_logic_vector(0 downto 0) := (others => 'X'); -- address
			simple_soma_0_m_synapse_waitrequest                  : out std_logic;                                       -- waitrequest
			simple_soma_0_m_synapse_read                         : in  std_logic                    := 'X';             -- read
			simple_soma_0_m_synapse_readdata                     : out std_logic_vector(7 downto 0);                    -- readdata
			simple_synapse_0_s_synapse_read                      : out std_logic;                                       -- read
			simple_synapse_0_s_synapse_readdata                  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- readdata
			simple_synapse_0_s_synapse_waitrequest               : in  std_logic                    := 'X'              -- waitrequest
		);
	end component test_mm_interconnect_1;

	component test_mm_interconnect_2 is
		port (
			clk_0_clk_clk                                        : in  std_logic                    := 'X';             -- clk
			simple_soma_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                    := 'X';             -- reset
			simple_soma_0_m_time_address                         : in  std_logic_vector(0 downto 0) := (others => 'X'); -- address
			simple_soma_0_m_time_waitrequest                     : out std_logic;                                       -- waitrequest
			simple_soma_0_m_time_read                            : in  std_logic                    := 'X';             -- read
			simple_soma_0_m_time_readdata                        : out std_logic_vector(7 downto 0);                    -- readdata
			simple_synapse_0_s_time_address                      : out std_logic_vector(7 downto 0);                    -- address
			simple_synapse_0_s_time_read                         : out std_logic;                                       -- read
			simple_synapse_0_s_time_readdata                     : in  std_logic_vector(7 downto 0) := (others => 'X'); -- readdata
			simple_synapse_0_s_time_waitrequest                  : in  std_logic                    := 'X'              -- waitrequest
		);
	end component test_mm_interconnect_2;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal simple_soma_0_m_spike_waitrequest                        : std_logic;                    -- mm_interconnect_0:simple_soma_0_m_spike_waitrequest -> simple_soma_0:m_spike_waitrequest
	signal simple_soma_0_m_spike_address                            : std_logic;                    -- simple_soma_0:m_spike_address -> mm_interconnect_0:simple_soma_0_m_spike_address
	signal simple_soma_0_m_spike_write                              : std_logic;                    -- simple_soma_0:avs_m_write_spike -> mm_interconnect_0:simple_soma_0_m_spike_write
	signal simple_soma_0_m_spike_writedata                          : std_logic_vector(7 downto 0); -- simple_soma_0:avs_m_writedata_spike_time -> mm_interconnect_0:simple_soma_0_m_spike_writedata
	signal mm_interconnect_0_simple_synapse_0_s_spike_waitrequest   : std_logic;                    -- simple_synapse_0:s_spike_waitrequest -> mm_interconnect_0:simple_synapse_0_s_spike_waitrequest
	signal mm_interconnect_0_simple_synapse_0_s_spike_write         : std_logic;                    -- mm_interconnect_0:simple_synapse_0_s_spike_write -> simple_synapse_0:avs_s_write_spike
	signal mm_interconnect_0_simple_synapse_0_s_spike_writedata     : std_logic_vector(7 downto 0); -- mm_interconnect_0:simple_synapse_0_s_spike_writedata -> simple_synapse_0:avs_s_writedata_spike_time
	signal simple_soma_0_m_synapse_readdata                         : std_logic_vector(7 downto 0); -- mm_interconnect_1:simple_soma_0_m_synapse_readdata -> simple_soma_0:avs_m_readdata_synapse
	signal simple_soma_0_m_synapse_waitrequest                      : std_logic;                    -- mm_interconnect_1:simple_soma_0_m_synapse_waitrequest -> simple_soma_0:m_synapse_waitrequest
	signal simple_soma_0_m_synapse_address                          : std_logic;                    -- simple_soma_0:avalon_master_1_address -> mm_interconnect_1:simple_soma_0_m_synapse_address
	signal simple_soma_0_m_synapse_read                             : std_logic;                    -- simple_soma_0:avs_m_read_synapse -> mm_interconnect_1:simple_soma_0_m_synapse_read
	signal mm_interconnect_1_simple_synapse_0_s_synapse_readdata    : std_logic_vector(7 downto 0); -- simple_synapse_0:avs_s_readdata_synapse -> mm_interconnect_1:simple_synapse_0_s_synapse_readdata
	signal mm_interconnect_1_simple_synapse_0_s_synapse_waitrequest : std_logic;                    -- simple_synapse_0:s_synapse_waitrequest -> mm_interconnect_1:simple_synapse_0_s_synapse_waitrequest
	signal mm_interconnect_1_simple_synapse_0_s_synapse_read        : std_logic;                    -- mm_interconnect_1:simple_synapse_0_s_synapse_read -> simple_synapse_0:avs_s_read_synapse
	signal simple_soma_0_m_time_waitrequest                         : std_logic;                    -- mm_interconnect_2:simple_soma_0_m_time_waitrequest -> simple_soma_0:avs_m_waitrequest
	signal simple_soma_0_m_time_readdata                            : std_logic_vector(7 downto 0); -- mm_interconnect_2:simple_soma_0_m_time_readdata -> simple_soma_0:avs_m_readdata_time
	signal simple_soma_0_m_time_address                             : std_logic;                    -- simple_soma_0:avs_m_address -> mm_interconnect_2:simple_soma_0_m_time_address
	signal simple_soma_0_m_time_read                                : std_logic;                    -- simple_soma_0:avs_m_read_time -> mm_interconnect_2:simple_soma_0_m_time_read
	signal mm_interconnect_2_simple_synapse_0_s_time_readdata       : std_logic_vector(7 downto 0); -- simple_synapse_0:avs_s_readdata_time -> mm_interconnect_2:simple_synapse_0_s_time_readdata
	signal mm_interconnect_2_simple_synapse_0_s_time_waitrequest    : std_logic;                    -- simple_synapse_0:avs_s_waitrequest -> mm_interconnect_2:simple_synapse_0_s_time_waitrequest
	signal mm_interconnect_2_simple_synapse_0_s_time_address        : std_logic_vector(7 downto 0); -- mm_interconnect_2:simple_synapse_0_s_time_address -> simple_synapse_0:avs_s_address
	signal mm_interconnect_2_simple_synapse_0_s_time_read           : std_logic;                    -- mm_interconnect_2:simple_synapse_0_s_time_read -> simple_synapse_0:avs_s_read_time
	signal rst_controller_reset_out_reset                           : std_logic;                    -- rst_controller:reset_out -> [mm_interconnect_0:simple_soma_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:simple_soma_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_2:simple_soma_0_reset_sink_reset_bridge_in_reset_reset, simple_soma_0:rst, simple_synapse_0:rst]
	signal reset_reset_n_ports_inv                                  : std_logic;                    -- reset_reset_n:inv -> rst_controller:reset_in0

begin

	simple_soma_0 : component simple_soma
		generic map (
			THRESHOLD  => 10,
			TIME_WIDTH => 8
		)
		port map (
			clk                        => clk_clk,                             --      clock.clk
			rst                        => rst_controller_reset_out_reset,      -- reset_sink.reset
			avalon_master_1_address    => simple_soma_0_m_synapse_address,     --  m_synapse.address
			avs_m_read_synapse         => simple_soma_0_m_synapse_read,        --           .read
			avs_m_readdata_synapse     => simple_soma_0_m_synapse_readdata,    --           .readdata
			m_synapse_waitrequest      => simple_soma_0_m_synapse_waitrequest, --           .waitrequest
			m_spike_address            => simple_soma_0_m_spike_address,       --    m_spike.address
			avs_m_write_spike          => simple_soma_0_m_spike_write,         --           .write
			avs_m_writedata_spike_time => simple_soma_0_m_spike_writedata,     --           .writedata
			m_spike_waitrequest        => simple_soma_0_m_spike_waitrequest,   --           .waitrequest
			avs_m_address              => simple_soma_0_m_time_address,        --     m_time.address
			avs_m_waitrequest          => simple_soma_0_m_time_waitrequest,    --           .waitrequest
			avs_m_read_time            => simple_soma_0_m_time_read,           --           .read
			avs_m_readdata_time        => simple_soma_0_m_time_readdata        --           .readdata
		);

	simple_synapse_0 : component simple_synapse
		generic map (
			THRESHOLD  => 10,
			TIME_WIDTH => 8
		)
		port map (
			clk                        => clk_clk,                                                  --      clock.clk
			rst                        => rst_controller_reset_out_reset,                           -- reset_sink.reset
			avs_s_read_synapse         => mm_interconnect_1_simple_synapse_0_s_synapse_read,        --  s_synapse.read
			avs_s_readdata_synapse     => mm_interconnect_1_simple_synapse_0_s_synapse_readdata,    --           .readdata
			s_synapse_waitrequest      => mm_interconnect_1_simple_synapse_0_s_synapse_waitrequest, --           .waitrequest
			avs_s_write_spike          => mm_interconnect_0_simple_synapse_0_s_spike_write,         --    s_spike.write
			avs_s_writedata_spike_time => mm_interconnect_0_simple_synapse_0_s_spike_writedata,     --           .writedata
			s_spike_waitrequest        => mm_interconnect_0_simple_synapse_0_s_spike_waitrequest,   --           .waitrequest
			avs_s_address              => mm_interconnect_2_simple_synapse_0_s_time_address,        --     s_time.address
			avs_s_waitrequest          => mm_interconnect_2_simple_synapse_0_s_time_waitrequest,    --           .waitrequest
			avs_s_read_time            => mm_interconnect_2_simple_synapse_0_s_time_read,           --           .read
			avs_s_readdata_time        => mm_interconnect_2_simple_synapse_0_s_time_readdata        --           .readdata
		);

	mm_interconnect_0 : component test_mm_interconnect_0
		port map (
			clk_0_clk_clk                                        => clk_clk,                                                --                                      clk_0_clk.clk
			simple_soma_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                         -- simple_soma_0_reset_sink_reset_bridge_in_reset.reset
			simple_soma_0_m_spike_address(0)                     => simple_soma_0_m_spike_address,                          --                          simple_soma_0_m_spike.address
			simple_soma_0_m_spike_waitrequest                    => simple_soma_0_m_spike_waitrequest,                      --                                               .waitrequest
			simple_soma_0_m_spike_write                          => simple_soma_0_m_spike_write,                            --                                               .write
			simple_soma_0_m_spike_writedata                      => simple_soma_0_m_spike_writedata,                        --                                               .writedata
			simple_synapse_0_s_spike_write                       => mm_interconnect_0_simple_synapse_0_s_spike_write,       --                       simple_synapse_0_s_spike.write
			simple_synapse_0_s_spike_writedata                   => mm_interconnect_0_simple_synapse_0_s_spike_writedata,   --                                               .writedata
			simple_synapse_0_s_spike_waitrequest                 => mm_interconnect_0_simple_synapse_0_s_spike_waitrequest  --                                               .waitrequest
		);

	mm_interconnect_1 : component test_mm_interconnect_1
		port map (
			clk_0_clk_clk                                        => clk_clk,                                                  --                                      clk_0_clk.clk
			simple_soma_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                           -- simple_soma_0_reset_sink_reset_bridge_in_reset.reset
			simple_soma_0_m_synapse_address(0)                   => simple_soma_0_m_synapse_address,                          --                        simple_soma_0_m_synapse.address
			simple_soma_0_m_synapse_waitrequest                  => simple_soma_0_m_synapse_waitrequest,                      --                                               .waitrequest
			simple_soma_0_m_synapse_read                         => simple_soma_0_m_synapse_read,                             --                                               .read
			simple_soma_0_m_synapse_readdata                     => simple_soma_0_m_synapse_readdata,                         --                                               .readdata
			simple_synapse_0_s_synapse_read                      => mm_interconnect_1_simple_synapse_0_s_synapse_read,        --                     simple_synapse_0_s_synapse.read
			simple_synapse_0_s_synapse_readdata                  => mm_interconnect_1_simple_synapse_0_s_synapse_readdata,    --                                               .readdata
			simple_synapse_0_s_synapse_waitrequest               => mm_interconnect_1_simple_synapse_0_s_synapse_waitrequest  --                                               .waitrequest
		);

	mm_interconnect_2 : component test_mm_interconnect_2
		port map (
			clk_0_clk_clk                                        => clk_clk,                                               --                                      clk_0_clk.clk
			simple_soma_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                        -- simple_soma_0_reset_sink_reset_bridge_in_reset.reset
			simple_soma_0_m_time_address(0)                      => simple_soma_0_m_time_address,                          --                           simple_soma_0_m_time.address
			simple_soma_0_m_time_waitrequest                     => simple_soma_0_m_time_waitrequest,                      --                                               .waitrequest
			simple_soma_0_m_time_read                            => simple_soma_0_m_time_read,                             --                                               .read
			simple_soma_0_m_time_readdata                        => simple_soma_0_m_time_readdata,                         --                                               .readdata
			simple_synapse_0_s_time_address                      => mm_interconnect_2_simple_synapse_0_s_time_address,     --                        simple_synapse_0_s_time.address
			simple_synapse_0_s_time_read                         => mm_interconnect_2_simple_synapse_0_s_time_read,        --                                               .read
			simple_synapse_0_s_time_readdata                     => mm_interconnect_2_simple_synapse_0_s_time_readdata,    --                                               .readdata
			simple_synapse_0_s_time_waitrequest                  => mm_interconnect_2_simple_synapse_0_s_time_waitrequest  --                                               .waitrequest
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

end architecture rtl; -- of test
