-- test.vhd

-- Generated using ACDS version 21.1 842

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity test is
	port (
		addr_master_0_data_in_condiut        : in  std_logic_vector(7 downto 0)  := (others => '0'); --        addr_master_0_data_in.condiut
		addr_master_0_dbg_data_in_conduit    : out std_logic_vector(7 downto 0);                     --    addr_master_0_dbg_data_in.conduit
		addr_master_0_dbg_input_en_conduit   : out std_logic;                                        --   addr_master_0_dbg_input_en.conduit
		addr_master_0_dbg_output_en_conduit  : out std_logic;                                        --  addr_master_0_dbg_output_en.conduit
		addr_master_0_dbg_write_data_conduit : out std_logic_vector(7 downto 0);                     -- addr_master_0_dbg_write_data.conduit
		addr_master_0_dbg_write_to_conduit   : out std_logic_vector(31 downto 0);                    --   addr_master_0_dbg_write_to.conduit
		addr_master_0_input_en_conduit       : in  std_logic                     := '0';             --       addr_master_0_input_en.conduit
		addr_master_0_output_en_conduit      : in  std_logic                     := '0';             --      addr_master_0_output_en.conduit
		addr_master_0_write_to_conduit       : in  std_logic_vector(31 downto 0) := (others => '0'); --       addr_master_0_write_to.conduit
		clk_clk                              : in  std_logic                     := '0';             --                          clk.clk
		reset_reset_n                        : in  std_logic                     := '0'              --                        reset.reset_n
	);
end entity test;

architecture rtl of test is
	component addr_master is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			avm_m0_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			avm_m0_write       : out std_logic;                                        -- write
			avm_m0_writedata   : out std_logic_vector(7 downto 0);                     -- writedata
			avm_m0_address     : out std_logic_vector(31 downto 0);                    -- address
			rst                : in  std_logic                     := 'X';             -- reset
			data_in            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- condiut
			input_en           : in  std_logic                     := 'X';             -- conduit
			write_to           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- conduit
			output_en          : in  std_logic                     := 'X';             -- conduit
			dbg_data_in        : out std_logic_vector(7 downto 0);                     -- conduit
			dbg_input_en       : out std_logic;                                        -- conduit
			dbg_write_to       : out std_logic_vector(31 downto 0);                    -- conduit
			dbg_output_en      : out std_logic;                                        -- conduit
			dbg_write_data     : out std_logic_vector(7 downto 0)                      -- conduit
		);
	end component addr_master;

	component altera_avalon_mm_slave_bfm is
		generic (
			AV_ADDRESS_W               : integer := 32;
			AV_SYMBOL_W                : integer := 8;
			AV_NUMSYMBOLS              : integer := 4;
			AV_BURSTCOUNT_W            : integer := 3;
			AV_READRESPONSE_W          : integer := 8;
			AV_WRITERESPONSE_W         : integer := 8;
			USE_READ                   : integer := 1;
			USE_WRITE                  : integer := 1;
			USE_ADDRESS                : integer := 1;
			USE_BYTE_ENABLE            : integer := 1;
			USE_BURSTCOUNT             : integer := 1;
			USE_READ_DATA              : integer := 1;
			USE_READ_DATA_VALID        : integer := 1;
			USE_WRITE_DATA             : integer := 1;
			USE_BEGIN_TRANSFER         : integer := 0;
			USE_BEGIN_BURST_TRANSFER   : integer := 0;
			USE_WAIT_REQUEST           : integer := 1;
			USE_TRANSACTIONID          : integer := 0;
			USE_WRITERESPONSE          : integer := 0;
			USE_READRESPONSE           : integer := 0;
			USE_CLKEN                  : integer := 0;
			AV_BURST_LINEWRAP          : integer := 1;
			AV_BURST_BNDR_ONLY         : integer := 1;
			AV_MAX_PENDING_READS       : integer := 1;
			AV_MAX_PENDING_WRITES      : integer := 0;
			AV_FIX_READ_LATENCY        : integer := 0;
			AV_READ_WAIT_TIME          : integer := 1;
			AV_WRITE_WAIT_TIME         : integer := 0;
			REGISTER_WAITREQUEST       : integer := 0;
			AV_REGISTERINCOMINGSIGNALS : integer := 0;
			VHDL_ID                    : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			avs_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_address              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			avs_waitrequest          : out std_logic;                                        -- waitrequest
			avs_write                : in  std_logic                     := 'X';             -- write
			avs_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_begintransfer        : in  std_logic                     := 'X';             -- begintransfer
			avs_beginbursttransfer   : in  std_logic                     := 'X';             -- beginbursttransfer
			avs_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			avs_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			avs_read                 : in  std_logic                     := 'X';             -- read
			avs_readdatavalid        : out std_logic;                                        -- readdatavalid
			avs_arbiterlock          : in  std_logic                     := 'X';             -- arbiterlock
			avs_lock                 : in  std_logic                     := 'X';             -- lock
			avs_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			avs_transactionid        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- transactionid
			avs_readid               : out std_logic_vector(7 downto 0);                     -- readid
			avs_writeid              : out std_logic_vector(7 downto 0);                     -- writeid
			avs_clken                : in  std_logic                     := 'X';             -- clken
			avs_response             : out std_logic_vector(1 downto 0);                     -- response
			avs_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			avs_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			avs_readresponse         : out std_logic_vector(7 downto 0);                     -- readresponse
			avs_writeresponse        : out std_logic_vector(7 downto 0)                      -- writeresponse
		);
	end component altera_avalon_mm_slave_bfm;

	component test_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                        : in  std_logic                     := 'X';             -- clk
			addr_master_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			addr_master_0_m0_address                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			addr_master_0_m0_waitrequest                         : out std_logic;                                        -- waitrequest
			addr_master_0_m0_write                               : in  std_logic                     := 'X';             -- write
			addr_master_0_m0_writedata                           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			mm_slave_bfm_0_s0_address                            : out std_logic_vector(15 downto 0);                    -- address
			mm_slave_bfm_0_s0_write                              : out std_logic;                                        -- write
			mm_slave_bfm_0_s0_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			mm_slave_bfm_0_s0_byteenable                         : out std_logic_vector(3 downto 0);                     -- byteenable
			mm_slave_bfm_0_s0_waitrequest                        : in  std_logic                     := 'X'              -- waitrequest
		);
	end component test_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal addr_master_0_m0_waitrequest                    : std_logic;                     -- mm_interconnect_0:addr_master_0_m0_waitrequest -> addr_master_0:avm_m0_waitrequest
	signal addr_master_0_m0_address                        : std_logic_vector(31 downto 0); -- addr_master_0:avm_m0_address -> mm_interconnect_0:addr_master_0_m0_address
	signal addr_master_0_m0_write                          : std_logic;                     -- addr_master_0:avm_m0_write -> mm_interconnect_0:addr_master_0_m0_write
	signal addr_master_0_m0_writedata                      : std_logic_vector(7 downto 0);  -- addr_master_0:avm_m0_writedata -> mm_interconnect_0:addr_master_0_m0_writedata
	signal mm_interconnect_0_mm_slave_bfm_0_s0_waitrequest : std_logic;                     -- mm_slave_bfm_0:avs_waitrequest -> mm_interconnect_0:mm_slave_bfm_0_s0_waitrequest
	signal mm_interconnect_0_mm_slave_bfm_0_s0_address     : std_logic_vector(15 downto 0); -- mm_interconnect_0:mm_slave_bfm_0_s0_address -> mm_slave_bfm_0:avs_address
	signal mm_interconnect_0_mm_slave_bfm_0_s0_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:mm_slave_bfm_0_s0_byteenable -> mm_slave_bfm_0:avs_byteenable
	signal mm_interconnect_0_mm_slave_bfm_0_s0_write       : std_logic;                     -- mm_interconnect_0:mm_slave_bfm_0_s0_write -> mm_slave_bfm_0:avs_write
	signal mm_interconnect_0_mm_slave_bfm_0_s0_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:mm_slave_bfm_0_s0_writedata -> mm_slave_bfm_0:avs_writedata
	signal rst_controller_reset_out_reset                  : std_logic;                     -- rst_controller:reset_out -> [addr_master_0:rst, mm_interconnect_0:addr_master_0_reset_sink_reset_bridge_in_reset_reset, mm_slave_bfm_0:reset]
	signal reset_reset_n_ports_inv                         : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0

begin

	addr_master_0 : component addr_master
		port map (
			clk                => clk_clk,                              --          clock.clk
			avm_m0_waitrequest => addr_master_0_m0_waitrequest,         --             m0.waitrequest
			avm_m0_write       => addr_master_0_m0_write,               --               .write
			avm_m0_writedata   => addr_master_0_m0_writedata,           --               .writedata
			avm_m0_address     => addr_master_0_m0_address,             --               .address
			rst                => rst_controller_reset_out_reset,       --     reset_sink.reset
			data_in            => addr_master_0_data_in_condiut,        --        data_in.condiut
			input_en           => addr_master_0_input_en_conduit,       --       input_en.conduit
			write_to           => addr_master_0_write_to_conduit,       --       write_to.conduit
			output_en          => addr_master_0_output_en_conduit,      --      output_en.conduit
			dbg_data_in        => addr_master_0_dbg_data_in_conduit,    --    dbg_data_in.conduit
			dbg_input_en       => addr_master_0_dbg_input_en_conduit,   --   dbg_input_en.conduit
			dbg_write_to       => addr_master_0_dbg_write_to_conduit,   --   dbg_write_to.conduit
			dbg_output_en      => addr_master_0_dbg_output_en_conduit,  --  dbg_output_en.conduit
			dbg_write_data     => addr_master_0_dbg_write_data_conduit  -- dbg_write_data.conduit
		);

	mm_slave_bfm_0 : component altera_avalon_mm_slave_bfm
		generic map (
			AV_ADDRESS_W               => 16,
			AV_SYMBOL_W                => 8,
			AV_NUMSYMBOLS              => 4,
			AV_BURSTCOUNT_W            => 3,
			AV_READRESPONSE_W          => 8,
			AV_WRITERESPONSE_W         => 8,
			USE_READ                   => 0,
			USE_WRITE                  => 1,
			USE_ADDRESS                => 1,
			USE_BYTE_ENABLE            => 1,
			USE_BURSTCOUNT             => 0,
			USE_READ_DATA              => 0,
			USE_READ_DATA_VALID        => 0,
			USE_WRITE_DATA             => 1,
			USE_BEGIN_TRANSFER         => 0,
			USE_BEGIN_BURST_TRANSFER   => 0,
			USE_WAIT_REQUEST           => 1,
			USE_TRANSACTIONID          => 0,
			USE_WRITERESPONSE          => 0,
			USE_READRESPONSE           => 0,
			USE_CLKEN                  => 0,
			AV_BURST_LINEWRAP          => 1,
			AV_BURST_BNDR_ONLY         => 1,
			AV_MAX_PENDING_READS       => 1,
			AV_MAX_PENDING_WRITES      => 0,
			AV_FIX_READ_LATENCY        => 0,
			AV_READ_WAIT_TIME          => 1,
			AV_WRITE_WAIT_TIME         => 0,
			REGISTER_WAITREQUEST       => 0,
			AV_REGISTERINCOMINGSIGNALS => 0,
			VHDL_ID                    => 0
		)
		port map (
			clk                      => clk_clk,                                         --       clk.clk
			reset                    => rst_controller_reset_out_reset,                  -- clk_reset.reset
			avs_writedata            => mm_interconnect_0_mm_slave_bfm_0_s0_writedata,   --        s0.writedata
			avs_address              => mm_interconnect_0_mm_slave_bfm_0_s0_address,     --          .address
			avs_waitrequest          => mm_interconnect_0_mm_slave_bfm_0_s0_waitrequest, --          .waitrequest
			avs_write                => mm_interconnect_0_mm_slave_bfm_0_s0_write,       --          .write
			avs_byteenable           => mm_interconnect_0_mm_slave_bfm_0_s0_byteenable,  --          .byteenable
			avs_begintransfer        => '0',                                             -- (terminated)
			avs_beginbursttransfer   => '0',                                             -- (terminated)
			avs_burstcount           => "001",                                           -- (terminated)
			avs_readdata             => open,                                            -- (terminated)
			avs_read                 => '0',                                             -- (terminated)
			avs_readdatavalid        => open,                                            -- (terminated)
			avs_arbiterlock          => '0',                                             -- (terminated)
			avs_lock                 => '0',                                             -- (terminated)
			avs_debugaccess          => '0',                                             -- (terminated)
			avs_transactionid        => "00000000",                                      -- (terminated)
			avs_readid               => open,                                            -- (terminated)
			avs_writeid              => open,                                            -- (terminated)
			avs_clken                => '1',                                             -- (terminated)
			avs_response             => open,                                            -- (terminated)
			avs_writeresponserequest => '0',                                             -- (terminated)
			avs_writeresponsevalid   => open,                                            -- (terminated)
			avs_readresponse         => open,                                            -- (terminated)
			avs_writeresponse        => open                                             -- (terminated)
		);

	mm_interconnect_0 : component test_mm_interconnect_0
		port map (
			clk_0_clk_clk                                        => clk_clk,                                         --                                      clk_0_clk.clk
			addr_master_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                  -- addr_master_0_reset_sink_reset_bridge_in_reset.reset
			addr_master_0_m0_address                             => addr_master_0_m0_address,                        --                               addr_master_0_m0.address
			addr_master_0_m0_waitrequest                         => addr_master_0_m0_waitrequest,                    --                                               .waitrequest
			addr_master_0_m0_write                               => addr_master_0_m0_write,                          --                                               .write
			addr_master_0_m0_writedata                           => addr_master_0_m0_writedata,                      --                                               .writedata
			mm_slave_bfm_0_s0_address                            => mm_interconnect_0_mm_slave_bfm_0_s0_address,     --                              mm_slave_bfm_0_s0.address
			mm_slave_bfm_0_s0_write                              => mm_interconnect_0_mm_slave_bfm_0_s0_write,       --                                               .write
			mm_slave_bfm_0_s0_writedata                          => mm_interconnect_0_mm_slave_bfm_0_s0_writedata,   --                                               .writedata
			mm_slave_bfm_0_s0_byteenable                         => mm_interconnect_0_mm_slave_bfm_0_s0_byteenable,  --                                               .byteenable
			mm_slave_bfm_0_s0_waitrequest                        => mm_interconnect_0_mm_slave_bfm_0_s0_waitrequest  --                                               .waitrequest
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

end architecture rtl; -- of test
