`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IOEnQI1AgEvONg23kl+qnHlK9OlmqlJzX0tPT8qeVEMisJEEtEc5YsVk4t900NVj
i96dZqUDun0uxw1SEEegxsoZbWMwzjHjD0QkRgVlGesawTz2cR/4XKZoslvFl+Wy
bQeQ+ve8n6MLV40JF6DNxM/1LM5l0H0X7DqOsUA5ABs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2848)
FdiQb0tX6AqxBXbxsbPu6kvP8/dLUth2wIowM6gaQZKnu+pi/yhFAEbEpp9AzaDO
evaWW3wfs589wCOh05fdsiYhtaZiUdzSQmQ4apdu091msecfeoRZnJaVfk1vCdXY
8ZLUI+e2sQ9TlbBxNgpdZPLdQ4MEkSHhDC2jYJ13Aj8XDC7DnZF3d1rAWhZtN3wX
v+0JbsrW9/izUCbrQ+q+dLOkH+NLlk+b1qBAICXY1Tx8UB2EEV3vVnrvK8attaHc
QnoZ30Gnc48etPo3UD41xNFjprgyRzD+a1yhEqUJkm0qchwWFVZXRYcZYRdMs1mM
xopbMcUJD/h1vvm6urgFZ8tQj43XFF+Q+qu7WVDtgfYg3h4gjUjJ66RIqgCkY719
wInSa/WWOwydsWbhaKG/JGxY9WJ8gEopLyV8vcVgj97hbqrPgb6gdkP0ZA9BrxJF
BuXE/rcHyyvBQIySFyM3FmC0Eck+//AQcUfybSnLkSQaJqha+3jovzEpeWsvUGFR
BehrcR6Dq8shglV3kC70KbpDSyfUnqufuAufoKdOg6h6/YadodjAxtS4drP9bcwI
nD0AJZ0dEHO+i5LSP+LsooeD6J5ETfuzD1Jroly9XXaGtWHWlv4A4egUXMycBUz+
VCQ81FfAC9ivdqHmGn0LQhKVI1BccwNIiWNzNA/pFc7N5/zb9h/40TdnDuWmgH7e
7Ns93DaZEvfluFfCIOsmuEZEY+5JqzwtnCHuSdSS7IvQXLi+SuBwftI4ErjJkBle
+5fVJgNqFhxQxcpaTXqtiCIFGlkUAXJMYfNgZAWIeCjQIyB+mB7Bo10am4jcOHyX
j2njkii45imJUPMf2AD4IdqFNgh2QTfpZ3dC8UHJ/RTzrJq0vRoGbSwwEPlxI0E+
OAHe4dpurTMLUx8/1krjnvEtquoP5pFeAAfFq3jMJot7MGC783V3wPb66jvh1fcs
pZPnBlpnU9aY+1WnVrXaoXdVZjHewfDYkFdnHU300SwaFZ3iwOffYBQq8TgqzwBd
8u08LbV2StuTEVmE8y/G/zfZimSLR/LlsqMxsVu9DgZMNXNhj5EVjlvpDqVPDBVH
EngQiiBc9xN9auRxGy9i4160ZSUpG7kY0HlyWHknvm58MpSUj7yjc/FyILxwItup
X14+d9oFyu9oq+xDoAQ/YUwoah5/6q87XMPEyVKaU5B1rgrYTu5pgLvfw1R95Fy8
SSRFUJtYCJGGZZ0L2bucVObOoSlLqt5mrf/tJHiJ9SvEc7YG8ZumAPuv7JwTzZYu
3xACfU+DmIsciz5etABRwvjr3p4wzVRaZtAHEUOmumhkk/yGVbuxhq/LhEXI8O7t
O+92m3Wb1A3HFxteAmHYT7yY5tTgMgycmtFlh2HHyYRnLY9VpnZna1igI0Y1UjXb
wCZvHGJ367dlBVEhZxwRYsCqZYkW0UE3CSY9/t4PeHeoasQ/e2oIwaetdLxLKmBL
bAL+lY6wFEq903ra+UMdzawfk5KjL68f+ZSz9F6+xHJ8MeT7iIeRc1mIIUjZGxqS
d+wld/FS3GSFvihrPA4PVoUpjlH1qBf/F8lJsPU7gQtO98BZ6ubaBPNXkJYcD4/0
jyg7zCJZzz82KQoXXWZFgapWDxu1ljzq0dewSnmJfPtU09GYjdLuXuXUynSmqsG8
lo9YoHaiQ14d7FMrkUXaASux+z+PKCe+N47ULuyF4oXMKKZofKCmttAlVCzdB328
GDlWypcnlfDUGL1tzlIHFD3QTIuxqXnDlrZFhvixHMJVYw3M6hauRAO7rM5cQSGP
e8h5SvRJvkPB/ZliC/qpDi8jdpOXcNPbn36sNJPS8W0b0zJQrHm76lK4o+cOSVdH
7IlvAg93/8EW66DcK3u6VvP4fzzBY7vfUVxeckbdn4GrttkTTVwm3LlooqIk2hRm
hGLss3ya68J0kVIr7xyDaEpYrVoRmjKSDC+Ymy5++bX0mOFzt2hMNWpvHGErQqNX
n4g3O5iGOMkEjr6nvVsgMQlIZQijqdVG5XK28S0NtP11aEjtYDLiKErVOfhIjGcJ
lkI3fV1Z3CUZC/dYh0fLPGKc+h6thd4dbkFRDojOfPYKTksIEfvgizcYhD6+fD6/
RejHChFpz5Hk7Ufa9A2b/hoe/JVAUJzejVpssP5LkC43/iK4b7zjFpMfaOpHtQiN
xoKbZOoBbHE9P1WHDSqaE5cP7WaKuzuk1dxGVdYpmyPfoCkYObUGAwGzs9pdaRq4
MiJMaOlEBhb//P6A2Ud8en8hJHCywI38++G1YP9nkj5g6TCEW7M/sfLR69+4tiUe
IeUp2awo4Ha2FBOSvI7/Xuu9sMav9Ik3UtUWS9yxgHBNfhcdThKRR4ODatct1ouh
W2SOnanLisRkiWnLUQko2LIJo0U/Fpj54wEpSXbTzzf3Mf6tFac1ZrNlmu/KN6xU
sluAnHa8OyXc+rQVOt7T6i3BOoiwgeud8J7qa59f727AmRhsCQ2i5QMThfrrQXWM
3N+yYAV7oQxiadNXSNgc47F8a9VflG5TuWCbnrELEZZwFjJ63609Se3sn98a3xoC
/M5dQYIwob09lGl960eR6ft/kWJVc4Lm5NvZi1OeMPSzHenr+ykoctABb26S4p7L
qxZVRO41xh7n29f2cQV3zL7Uy09XFLWQuYUVpPYA5kI0UWl24Mhf4Nk+D+9B/mrV
Xe3qm8VEt3W7ue2gJ4HAS0bCOQ023xkFLchvtvk+FOc13OGDeF02771GUBLUcAkV
+KYPnoqPJBnPu/EvfuK/CYntSY8Yyayw/Zfv8of+yOYfGjICPSm5l3I1JpcjiSN4
v6wR6zVOeVozMAjaH0d8M5VZb0zy9DpCJ3V8LeZnpncWL+aAzVqGX5gnCcgyn616
vc7mi1iGg2ldwdMrdjBtwlrUHZT40J91SYR/pqzOZ/kdXgwiU5SC1/SEWxTvwWrH
UuUlWUe8sLgG48NgYtgBGWJC+NGpExIMBi7vMgf28NPuXizIntjG9fGmcFp8bjQ+
giZsoHXLN7rOcjC7jD/+oICoWM2+CPg+mjaE8cSo2BGmKt4PVVJ6LTPHgLaQXjn5
btw18snnhKKVd/VU9Wmaw4mzSLXFwTHB3dTN7UoU+fKpBY9861j3koUQ269YcOWk
r3AdUfMFpiScyzk/1/lS2jH1DSYsWzSovf4x2RPFu2AObBMVIjFUAu1vzxJoDktE
AGZd83jow0LgKnQ1RMk9pHCd8770bnsWsMdTIHFgHLrB98wdXqH/Z6ONyEprNgiT
w/Hm1RIY0xLiUdyj16h0HnmVp6AWdaazfE3o2Ub6y6x4RZZ2xS7aBbSs3quS4ZrO
c4PAcZI7BgfXwGgwZZjCqOmyr7cgHeEciaudq3+uqYxKJht/AtVJzgQaTw1cci6x
mimmZtIONSp6vYFnS47AO2tp4PqpWCLUjmwVstt1hkCEoYko/CTbn0CdCBTIkbay
j+u5gZyhctVzbu4bYLQfS+U91WLsWUCSSIfhKlZsFjkeDIMiDBWPKDyPPcfFuSWK
N+H+C8HhkTw7m7ptnwaD7PByYHCFLabJVMCl/Fhj2AVxq03AZlL4x9TpB4gGdQdQ
TdKpam73SZ1Av+8Lc8DW13xu1hrlcm7aiJ/v2t6zz+gC0S6znPiWmihDkMFLEyj9
3hHiiYL4Oh4HPbqBmx2Sd6pdJT6zeElljU5f0hDkD4FSCWnu6yJM8oAM/Kev96rW
bCakm/xYQVnYVkob4ZfNMZpM9qHrDDaYgORDauKlWbD+I3ZNgFzwRysH8SQznYCZ
/iNKBr0QDKFnV3FMPk+mfA==
`pragma protect end_protected
