`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gmdNnLoW17IugU7VL1XkanMjpjXyzdCqDePZs+ChoFiZAcp76ntStiY1ftqILZHs
yZeUo8FbeCahE2dRfjBTwswWCXM0jc18AQpZxRR1NVSmyc6Se6ej2SQDuE3GAhqg
aus7cHKP55KVSGnC/5js2HDE2vH6gzHo4PdI2KX2bPc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29344)
vmYB4XOZbCkAXiYeWp3CSdqG8f1scxunKeH5fhllS2IxBKGriNqfyGFB9wX0pUU7
AoZruIk+xxOQQNZhjOtFsKUGJrdrRQi1YV9U16ZONhDjzUf2LNfnIckFyWXz5PfD
EVvpqcY67n7pzB2AIsQC8Cc59zqKuJ31yJMbltyjtZqtbqFoz2Pjfh+/1e9Ctgp3
+/rcAJF3gK9CqMevzdaKX7pb6HLb4cAHif4dMmH1a9IFXcdm2yv7k6TxM6zhOi+u
2P/zStpFBdDMShVR55sdrWDabwJVdpwwa9+Rz52OUIHGioVBoE0Huy4tE6lBu4ca
iiKXFppk5rm4hn79BNuWBL/9Pb8eJOzdDBZdn5tJaiRaFFBT56UDR0p91MEOHBND
Xc0rQsTao+fSV/po4FQEcZ6cb7MdZG+6CObq5atbDnRj6f/xk/mQimjQw3pY4YoY
LIL3cTvkL+T2g4PZa3KqDkla2hATiT2QAWzKpXdYTaiBSdwk254XBCdYNnu4rLDs
nMmjBu1h52c0P0et1pIiUW+hX6KRnXJvrYRbtLIBtWlimF8shRBQ5uEKZGrh9XNh
exl0YULI6dGmftYPo/skj7GAjqanqwB/1MbQZla5ASxwMyCIGeoZNdl81ZuL5mZH
6KGLVZWRiSM+5HfV11d6N9zL/NGnhY2TDWiJpEwGQx6jAAMgnf8iWtEuEd/aoUzT
GvMIBMxGn3K6oed7mna9so5CmhiWHI/h6OhI+3K3gDuAdC0mOptvImpRRec2+1xt
JkMm92QVePFgmePZBCYrFQRjeXiv+O/ID+vRw30LOu5ztt1W41Yil3S0fYl7hvb7
eabKKJU5rCnY4QRa1uoABgxyEsmOkzZ/pYuvjCELCdQ0CMcFsSKGdmNf8u4Pkw37
q7mDvrfzdliwEf8YpOVf/DXzrUMwXla9eQw+UsrzqZTZS9gR9AQ0akR+sYefgPjA
XCW2OTwucx5RrrnCN5BCXfvYBRuueW/Fg9v422Cyve4wb994fQ5uKkXzoLNBfojl
J5OTQXo8CCwoVlod/jDdcugbzJ6J6FnhamUjSRWh/wt4mLCvuUDf9pU7Lh/SahZ7
OS8ZJywN12qBkVjfT3R1pxg5gCkIbilmAEBKWSIu/g4F1HLk94NVclFTl61wF36/
UpI68TwDA+Jkhq2dAd2jkaEH5tl/kwLf34joxdNKlITxd1XERQxUku3StLiZtuKm
u8aa3967VtIHaUvu31Q5XCztakcUDqBiayg97AtKriLbu5Gz3HGJx+N+y1MCdNhS
fIRdQYtrBA6X4vneqcTcih+3Ig8o/6WU29HriXnINNYiv/I+oEWyMFXtHJSmthT4
EihnJE4ySmtHbxfAOEtc/zxWC0B09DlX2zIEKkeBYOfdm6yBi8l0cGV7omyuKz86
RXISSVOn/t1Ub9xk0zqV+xnG4+VSfjhkkpr9thlgdUTzZWS2OBQ8VuQ73tYDg3bI
hkW5C9FOveIvEZn2lYwoLgZelYuTYfedSrhCe/fOBYtXWdCJBGShRnCMBmjyO15U
cvFJfC3nW86Mb8qb6hBbK66VtrdXlgSQAWR0jTGufkxeuBswGLQe2VlIriOAfMl0
TPYEFD/4psqy+1Z1tPb2x+4vS/VS44Nfb5KUiBrcfTqmH4hp5VAvGm/Wk43FaXvf
6akUwMTQzue8Jo7k8+8LMn2MBmt67GMXhjwuXlFV+J9wJCYODR6AnCPJM9VNbZus
9xOVzvw/6hJJx15oa43DWpal5LsjlisacydrwQsI+Z6cU7LI7gL9ZimfNXEipEUp
8vLMjW3szXH98xjuT11c0EXBq80r/itjaILWaeIYNyG8PYiiFb7Edm4f3C51A3R/
FE1eKxxTHld/0N3pVWmKUyeuCbVd39WJwiT7vlqGvQlkSzZeECbh27QqaQpRv3Qy
pa6Bq+QuQBgyPw1ssJ6Lbr7B04qTC7/8bcMciRpWsqiZKwhfdGvlgIKJXsZOXkz+
NgltW82Ge40VJfCm1icjXygXfgvd1WQ8tfM7WNmB2qNoGh9GDnTn9NF2qa6SLIcO
rmjGla81/ROa1bqE9c6EZOk6wKy5q/nt0SQWicDnKeLXfzt8/ux903IBWg+zyk7a
Zzhcp3Aqxzg1KJqIxYYclWIBQOhs6+g8QimwDfJafwngkQutL11BV5hnOi8Bn0F/
12rlMuD6oNk456v1HjwuDe8BZI1Rx9JwPpPVhWCifpo+4RCu6kv3lyRw7Ct01Fz4
up2c+maEtbgHaufZAdnLo6gK4FockKgLkY95tnzI9l3KprzU9Tx+/Oeamjoe9aL5
kB4A/FtwoilPTxpMp9gWJhGQ8eTsUNI+eP2q8bTGMdZCbEh8+R86Qm9enheGjwJI
j/q2mlE/U4ow6B56Nwf9v9SSFYkC3hSZ5y4R6H0qjLkgicBaKL0+K5usgZS8EXjj
S5AoXGexbU8yf5xegDbjRpOmjozzIbGnpiA9liKqUCNi1Y9dFcnkh3XpbdlYAiUT
PeIlY0zsViaIsKK2UlHfrbVMqOqP9ejNH6EaOWu6zqxzIdVIWd8KDaMtXvKVvT7m
WxVX0f55KWcqLg7f5M0JXnZGqAbGj5SyoLlYel7WQh8gzN3f071hrNmgmS+a8QDj
G31TURG5l6PK71WJR+TxhxQuuezS+qZ24eyzMb0Y3+jh1xyoMqOdYkhWBTrLhwPc
0/7Cs0/DoK48Nl37ru/RYLXLaRTFaBc+bIQ2JBKEzs3VWHp4bkFRBE88P7J7c8yY
nSXu6l9hT+9NXAMguz25L3Ng5fRu88uey1FeD+XqrY0a8zrcQuhnlERUy8wLhzk/
YiracqXOO/sKNgNnEc04IfuDi/QmHtLSdbnQz+VamehMTMDlZ1rZiVB2sVDIigzX
ghVh2sKpgKNt2huPG5x1ToA/9EMwf/TZYL27ES7pnK68Q3sTzon5/ZkmdFwVUnJc
KodkIzePnL8vd9L8J2HSD3PB9XfINnu8HXd8lWX2E3exR9dD6827LT1N5/0LS+ML
yhO8Vlnc83EqLhuKGz9w/gwOxif7yVP72cHo8lKGf27jhp//0uPrRSG1rwdvieFQ
r5n7IuLTlFv3Rs50BG1W47rVEp2uzr08nJaBfBO9v6OAJEntErw51ALt28vtOLym
6gHeKjVHCZmcZQsChjTPExyPx134jIosJ+JyLsQWnyfX3i8U0NGzFdYFq2ft/Doh
PdiQTU0/rBQi9QjaIjhZm21h/0wc+JePjgi4y5Q71Le4mqD3kutGgcYmQz8NBezs
LtQe5n1yh9/F1oq30b1YKRIQoPhJnmMJYRd4YCPYOrfPvCTCqEYcEWEK4QL8/7rK
rUfRd8DJYVkao7ENppWQhP4OxQ06MEcWhHj9F5JpD8KfJa0aoan431bdNhHUBhE7
TbJI4VvCiUq0EOisBMm1Qr+PWluvFW00xqlciBxTK6EFQIxkAxa4yUs8w86uwWGg
MKLFxIog+aT8zN9whEtHCUaJmQd9CvRApO2z1bAmjaSpOfCcTbA7PLvG/AM0mGSh
PPHezh4HYe6+j8/bEwV+M8h1Zb5qcB5dkJECziu6VZ1c2iI2961KqC/iyhogZgJi
jI9qX/hD+BPMJ/lriwcMP6lkOsAbo2HKgGTq2azHxH+MqmpFUv5XqrLTOb/6561z
eL14/ft6TNLhCwMHKGuM71XAsjtRmOKPQGm4Mns+eG+36kBBAf7OtEoFb48cHjxt
x/pPfd5wK0ASUxiiR4hj4JwvSDlHVGGH2TsUZGj8zxAp8lAxSqHl/gZASVaBeM5r
Puo2yWgUk2nd4uWyuB7vZDmfX0DZbEREz3LH8IAx+QSm3xjoS88Xb524QGIUqt+9
I4ygLZZ40RWvZdX/qnPdagRn17fvyYQC4+JcNJwWF7YbsQPrwEKO50s4t7jA5Grn
5ltOrNq4Gtf98tX52rksr4jAj6kXbZaN+9OEh6+opZAHczCJIbsFVKt4fwTaGRSG
lVNWFHP3ogGAav0qp1DKUGAcyVfoTk/khVTBu0m8cTTxn7MPhfq/pfXWCPo6oAFv
XE5hm3QzxpdooSh59BRFShOwwryezEtHuxxSu0ZZ/KuvKGgplSq7jYdf/6ZUS7CQ
AU6F4tKvKUW8KzUai7ubYtH73knQ+Zio39EIlh8KM0n4hrr5XlpH9OPN4JY0APFD
ayS0oHiq6ReMT3Qql18kA3yIou5BbdDEXPwbqkrLvIEHLmN9lPTOmntX4EcuKI80
ofYeY1OmMt/y34h5BqKwhjJaAYwPvayrw2gL2YNtU0zhmCJUvm+yyQsXVci3301M
7mpg6kAWOR8X1jcRKhrZiU6CXzjmmv+ZpCdNtLanwoZCog0R/J2ozw8alwfVlXwC
dhLRvUOE9FjdBscUs/tQ30QbxKXYlm15YN8/Sx3SLxFNtHYtYC0D2OZ919rCZSMl
7HaG41q9oKCJX6ckDjixvP/KUQ0k8p8X2MmNDxtY9SsMozSSK9tkfpZ4eQomPxLd
bqlgJl4DXWOJMwwBvASxGhUK3S/R5KDlSFomDbdVB/Z9mMf/GEnWq4FjrtOZ/xnb
+bPPF/YeO8Ikx3gOOknxVclzTRQjXtHr9CMNpJQfKH6C8FrXuywma5oELoJ6e4/u
1s3ej7d2ilEIYZdv/Z29tEIi+lp7PVpcm3TJk1zoXaCrGRQHCGpWhbLtjd55N47h
OzYiYLkTk+DARdmWn4gH0uXAr2ChS8j4N2JeLbBz0CCzAsS6aD8vnOWxmUtrllpP
MIWX1vYSnDIMsKrfGiFqayClvYXOGdJrcAYHTc8jgsvEsLiStmVV31K7ti2NUcrG
F0bnYr8b8937Wzs1zmEOQUL7HYU735LPkxqFyAVTKhwegITFEHLbA3+ogIFzQdev
IoP92pInWa1N/84KVLwy0cPHKUe5C0FI0tBpawjl2vw/yKLAL1PGaML6lOvplfXx
eUULCIjlo4mKYIVqSKmWRNMeW6yvjVYzrh+OOvv3P2lEJz5BrWX4nvawnwvIWpBS
gFAL7pnQRNPmziitbDt4flfzkQ2yyoPgGzmVXd2b5m+BVCiwfAzBq+d8miHi9ooI
WbI21+5tS5/omKoPiGGR0KZGlb2aapVpLlLvndPQ3JKgAmWvgMlB65bNhtTHH/H5
/m04fHjAIEh5T/ZNMoqsT8jFbnzgC0XMiUirz5KJI/p2QiKSdzoT49hzymJM5AEa
gB5/KPe01PfE4V4vK5hmQWQNRyBXeQU5D51SueTF3izDJxXiI9xQnXod889G6mjk
phOvLd/xWncd4z0wI+xAhQQE104utzMmmQXBQi2O3gO/rCIJtI74/pxJSeiDSPTa
WcrEDxXymJRvSENnejBf4TClT7lJ1FAAxxA4Pt1hxafIEdvcZLN17ZMQB7P8YI2b
M4HdnESqd5G+NBlgtLK4dIGd9+a1nt4vBcwssj9lviGiancZR288XEmhzonotAYQ
WdQ/0JDgC13AaoFSldmqXHDgIWQDiLsQ1VqOL6HQzkGCe0fLVbZzMnt5+N1Nb5iR
D/l+CJoyE/+ywuSl8IkUvkxaOCjEGcyHeqRuDUgJmoWXk0ONhhKsS87eyfvwedk+
F+x+xLMgKN1+s+3lOHnzHaFK6pod1J9b9d7Eqpucn438GIsRjLHtjGK0Ruqf9F9G
FzgWY8KrCfBeSORfi7qg7cbwi5bADlJR+3KeNzlh4TygI008M4YAPW7L+NESx+fG
jcIRRL3EP88TOYPLEZTHSdRhJrmwJ/evj4w2hdp3jGcqw9A1b+dDccEK3F2eL3KP
9auGdwPdiy8PrD7EP+U/CybwvA+s+jh0tsRZYVIJjn6Ylb8sCk1/ooaTmm0NsjYK
IybicCJEO/MVhWMShqO8aDUkmfFPDcy+ROEDlGfW82SV2PdCl/YqqNulsV3Nx51r
ZP5odBYEgx768bfeCnEoF1SzLlpzASNEUH1QxxY4smlCB9L3WjoEa/idpUVbFnbx
l4RtKkOmTq+/mC/G4449wMS1L8H5Iet+TmicV615oJlXdXvz8UqpRyut0Ok5yspU
PVhJveralowWHcA3fxXK45tIB2V6jgxzDz4UGjIAUz1DZfwCa9vVIi/mFQJlwZus
VcJhVXfvJy3Gk5snvXUY1D8laVSgykxgl0NTuCGvWxKWla9bPJIroF8DeFTZ65Yu
t8b7WQKvC5MgjrxDwnn4PBc1nm/TZ2aA2lWMV+mntlOA52LuqL39KPje6P19V1MY
5DziXu9VJAKoizLUthbuiP2nSHHzysFDQdvi/k6zcg0HlwQA8IH9qBNux9YYuvIq
VJrUNSpinr9CTBR/99SlPqYK30IToTy3J2VMc9+NdtI6vW2JhTou14NpMzkip+nZ
e1NT+N1OJCaqtLvG4z9KdXNOaREqjuLNGU7p34OsJThrOIBKuLOqKIgZMFD53Xma
L8OH7ofXjlhoy2JL8otktgKeKhvzNSgS3QK7j5TNqNMWw6VvoSsKxBHJejAqWpzd
+HrKr1J1qkJEPb5cTafWc7F3jKgjiPX5vAOctflrk8wRwXivNUQ3GybOvIqa8NFW
LJwwzGvv+6a5WA9zEHmbvGijzHJAJa7HgYnHhhLxKc6ldkS6Xen79hsd0Ksvgaw6
ZPjK1X/21HVpdbAuZsMd582KNPtngjtFdlFaF0X82OoCjmt+namY36Viqacjmwd3
VUXZPFwVtaFDyhby0ir/U7NOnupvIfYJQ0KxrZ893lJlJEwm9uj8jye5XkFdVk84
fgYfrCVY6fE/rUjZ4h/EDU2hzgDthbkJykivndN//WclyDJRzoq91QkLmZ8yFydz
e3nJwUImyirqVRfmjElh5TCVoKxDef/Hn0XuobjvznWjEIu9Lx9ANVn9nSm54PZg
UF261DG+g/ILEvGKGTqL/UOfv+YAI+3LfwKTrNsWx88hPhBIlMxEAJUu1xdg7tl/
mAJvIbbLDQ+QONpvzGdlPfnOEAX6OT/R4iq36UU7n9yvFvLB9R131Lokcaz8yitv
r/ycxpnb64j/hzXg7/44QfGjSumHmPCGrVa+7f0vQTgeJGqR32pXwyd7R8BeocUf
ZjvowBRvvZAw7qIY+hYyzpef+JqFm7cPHPTlfcHT6fz9ocw3+4/CT+36HwN+Idll
uNs9XABGEvNbyYWAelKUm5drPzGK5jZ8dy/LkKF2m3r2FRojYCNa/xFP5b2rkTuP
PSOM63SU5eDbmZc28s+4SMZ29tst8iYFJgM4SbdluQT7a7ehE45bI0KBAfvceWwn
/LPDq6tLFn+HY3AKfPW4L5j+uMbElUEc7YnU6RBgcYpNYD8e8tABspZHN25CLKtA
3uW9CYcZCH/uMZ+4FJhXLZ67ETeNkxBctqRc6QASEmFt/tXehrQudMBS/57+6qUG
t+dCCKKDqLQCoF8/0eMUdEFYVO63uiC//pm0ZfkMxTke5C3duYaBkCBcnPy+TkA+
O/MYAqhaBrU7mIFrGZgJi5uUOI6Vtj/UwiJNX2HZVB8znFQLmmlPpV30h/lQpu29
VTytBZJ+TU68EV9oxyChCpy6IFRn57tWP5jWQkKNfPAt9gQEdYW1+6R+JuhZ8Css
6MGWJodT3odsDWdzfUmXCnIu+ToJ6s5Oz/ifcMk3pqQxcNi2mmGCwARSs6Npmv2H
2DmZxM43PVLgsyZ34qNMmI6pJni8I3Q8ZAFHPCOnBaJ29ldsMNoyKGXh2Tyg+yjF
8RWynjfUscG8VL+0PyjoIB3MUxLTIY/BxXwGU96MCVmZ/n/nPk/US/1fL2Z+Cny2
iVQVWEk3Eu6YLxqMtHe+Wss3EyHC9G8X/uSEYm/8rSjX1kQY2hmBaldVjCOhp2fr
uXajaAKwcgRVkOL1x8/JFcM3D1YXSKsQN/17OkOI/4XF536avV8KyKKehbb/ZLzj
QrLWi03bOQN42LY4JzDs4RcbdWZmU+XM0GJlBFyM15jRpGopNVnq9zxKQeWVTqRA
n/rvYx8s1dh6DSQA0TFsS1YA7HYvj2XI8DVGGw+4Y2cFj4HU+5XWiTB1Ut676pm9
zMVhoswGvbnIeKPOc7G/5jb87AqxXjkrKO0KCrUc5XWMHf4NhM0WRrhvH+GOrPUA
MAuP6wxEXa/k4fXJK7mbLJBp7TxWQoRjRye0lZ+8va8eRb54j8eUWNU7qglan7wj
9hBWH3Wb7OTjzyuQtqOleMnDx308ZVg+Xwy0E98B6KN1baTCMnH2QBfn6JFzoAzM
m5Uzqli2qf30bRbTqZJpEyCSVcCCWZmqT/x6Mh4nPj3TmezE2Wrj5QiG8VjfJ0Jt
EjsGE+9akzU9WaClo31qNHpRdMMyWgNWJQ2E4dH84fHwydUCGBZ3NOIZaUh9uq9C
3eQLWSwO/qPzy2gZETiv98W2aFWNfqVZ5ax3pwuk9GPecHE4eussPRaYvS1874TN
kz2p6RFlzVEVvnFRqmVWPffeItIxlXIVhtPx+8aq6p3fjtDUvAfgKhdd5OmA1a49
U+zlU/keNZaw9gdaBARGxET00OgZ8XkSVaUatN5/qzbxVIck14B5AG0K6WEb2yaB
Aad17P7FKpZlPibp6Dc7cofnIM5DeApdBLrJPw1UpgtjpKsPMH8/RavQBRxyEXEW
vVwRV7SheTh8B4WpxU19YsUlvmOxwJrDWVaRpqNXyXdnMRBHNWArimYgi/Zka0I0
pZ/fFbm9T3eoJFEGOGULkx0Kp3j+L1+tt/6PkE0SLXO4fcMEyAcMKqIVS0YZymCG
FUeq4+uF6PYtFORUi1tO+Cg71SS8lmKMlwG3CBROfbia7mlXztv2wOyTtZf9xql9
Na4Jy1s1/jNnT+zrHkxlTj5ROlpWaetMZufXVOh0r+aDWzdDmG9NJq9V22jwsdxs
My31RUQBVDLqyl4JiKUWOGAklxRF5eWR+FWjQ9seAleHWddnfB5d39e+M6VHrtQC
VfJQZCvZ1yA4E+i4uCJDYgq6FqeHdt7q81wp+ZsJEoclDUoXZS8noKiNr+dFK6ac
rd1xayTBOYjbEnvjL2a+HVzvLpNiG5GVttAx06g+DoZ1lnRnkCbJKlYWwx6wesQK
tLzXdE8iqRKkWhbdMzSHnelebMiUUsybqKm3awnRZcH3KvgVB3wJVuK1z0JRHL/V
R4iIcSQ6f957Cm4ty1Px4s/yFQGTnCp51k9zRuiTtQyfy5HnYt6npt4mJ83IaCTg
jOnVy+sDuhZ4Z/ve6N+8+8qaDeriLVbmKx3BZzALwlQTA056qL43a11OLZpzxi/D
EPKXtUM5A493PAwXvLudfkd6SYxJta1qxsC7FRVtQ0RPCsDJ4hwNfJQC6YiVTze8
EWCO0WIp6PG7R24pe85OpQofVRIo5Q4YPPavl33/EDVYSYld9mk5bXb4h9Z9qNsE
7rvugUiA9xhwgz4rsOMArYvUMjSTK+NKAOULKuLG459UkXWoVuZAuVxM+qgA0n3T
buAIdQwUQjGEg2ebfWIac4bSx3IisEyuAsEV5gwrbleDARy6NeHoP64BwvHLued4
/YwgicV+eJFF2vkxxJFJKtIprP0AsKhCCJdM06wGEGj+VLJHmea5b2oOb7Sn8drn
RsS6okYAwsMePEcF41CEtCav9dKx8DSA0jHMY/O/GktwXFalJcBhJ2EvsXNNcg5t
KhGaQFLWkL8/GB1xrQLKPwEOm8PHhuu2/8NZpYwbS+lM4+mZcFpF4WaxAXnNldUf
f+7wB1npWtCeVGeUtB/8pIsvhx1thl9K/PTr01+c+e+68JMVNqSC3fFCof9nF7M7
3qZItrRIOJo7o5DER3MnuoWrmUuqDj8H6m9XZ8pcoMM9WWc1LkXmLCagvAU9DcJS
JSM1UU4xAbOdeKqcOimxpjiawuCRpq4SJnd5Q0pSLQgimLXGIelliEmSPwP6Brwo
CSIiv4SasGdPKTuBB7LePGh/LEERV5NEDgPFpvddYpNQUp8iANEHwZ9l5Qk3rZ0u
XHOAtLzZTDKGKtY2Pr71w34LX6zUxzW+A5ylSEZbDYSvd8Ka71AGcdWgFDsnGAJL
kvhM+o7542sYd61lXVj1KNMMHZ09ewcOFP2/xpnCb+fNMF7pODy4Xjk+V7jJ7+ZH
8x519FqyAKXL/6IDzQX7FQyVqMhWa+9ax4rMVx9sd560xtXzvmxcfjb6hWV3TOct
qkNIXsbTNZ75HmLwRnI06g2neajMrqGId45gqSUJbMToUoDRoWNKpOlrvstx2jzE
dp+xGqR1SHdwU4UIksUEKYskbKp4XD/8davLw8ay8rw1Wy38nBGDkFepslt3WeSO
EIrbXOk5TTqOJo9c6wpSzv1IiDEjHO2Pa+MhMVlZM0Vx+hgaDvryfotdb3mEw6EY
4tLhZ5U2U9YWG4eFyQ323TFGJEtTzpCVU0V5QZ8Nvr9gvVIiTEzTPDC/NWOw4Gwe
310ekk9oUyD3hjU99d4PZsaNAETj+aouywB7Uj8/taBjNJgg8paGe7C/mHS3jvoh
OWSHiqAI1F+yE7fwsCE2YyDe/uBoawP0IZ8j1HSq1GYssjDLWkg4J9bKMwHfvoCm
nyI/EhDNRHXO6dKndZoxZpwFFM54k2vGJHnc6bemoHsS/bPyeKaDuE5BSsQQs2/g
aISsOnr67U/iyW5GtFwCn+1gBZsmp2e6xO4CUvgR+iU3T+hYQZ3W7X2uUhaXsjvw
yQUu7TpceutBdbRlpHO2onsy92YFC9DeeKg+8Ut7nDolY9dUIm7r02YSM6lmkQIb
xQKIXivMmL63ufSvX+0sbxWIFSPrYVoAzGTfI1UnU99R0Cgk5sAdI79MHn/sjtOT
Rl00NYWjxwqmigu2aubXsOAJAALoIYCYkDzbNz2Lq3Xb/yZQDWRaX0YpoegS781U
swPk2TrxyDhx7+eSC3dTSxNfl3JbFgAqE7XX0wRlu17t7s6Y+vA+soZWREWfsfiS
7/t7YwEmqv/sesAF5TByf343AKafGc/VlIs3Vkxai+z8QxirxcDlGDS/D+hOR+w7
rCDPI4YgDz/BWFFHQzn8TF24I0H1Z3OsgAXSAGl5IVKQ8z3LVDLQBW867SRFwbZN
1AT6uVV7sP4ktOlXXeOss28Xi9Zpz9JBJAeQ+f6m6WebRTL8VP87/OuBp0nbg3gn
176STcTM0MehqQpTnSkTGa5kKkYFMrRAWCtCNsWUrhXouzS2wfE9UPabtip8tCii
llqj6anpFx98F2jN3oCJ9TrxhjGEKEaLYZf1TTne71BziequapliLWqnrCweZvjw
PEGzMn7u1xCVYMngAPaePEGFkwIwza0hPdgN44GFH6wsszB4yBSs5FCMWUcL52an
iOVQQxr1m4cPeZELe3fXmIrbA5fHHUECEK5djGBmzNbgo6/uDdEqU8byjTvOy/bk
4E3t0ubV+RP8DbaLJOFd5ED0lns9ORXt3bWFH6GAR5oEwX2Rqw9HZfu0zonaqcJ+
SHfRc57xb+xzC0gj5jkyMZ0wDKQSrChXLUo41ae2MaGF8QdCBtkpIydI8yO4OYne
ZnjOTCGyq63dSSY62ypgUhETGQtKCXywPcpQDi5I8zIELQ/FNOIwCRpEZ4mGQpHR
XLUIBeCO5Awg9fSR1kfEnMy+lIe462B5+vMDCLRGrLkn1BEK6NaPbIqxvQ+GFulB
MftMtgBN1MPIgXysgF5EL9zaGYoi4Qo4reqKz/wz8V5xPqhA1DQMsRuJ55Ee89/Q
7/HWoDXH+/S+fzPJiggPjH6If+okT9jmQeDv8LEB/R72+QPLXysH6ihpbs1bBh8j
fCZaiTBNCU7Iv27XKfMC5QnMYhNrSE980FgRulJAooawUFyCKR6Wt0X49XHb/2rJ
cF8aAOcWk2HsbOq/UKg1SeRyisKaD9nEW9mTX/SM/vwng3mbXalt96fBavaihpga
dgmaihGSy5v5qHQSXjU76/PwW1roBvUnfN4DoUuupEf8AQq1WJ77NlaNv6NFUNAf
NYxXBhcYe12Gm4nJ3H+U8cFTRsHdNfHvoKawCwuwVMDVArTeHBzeLJd+8ogwMfmK
NYCd0+HIwahqkjUWVD7RFAZXIJIjVpD6bAtGjHjjAdBoLUlnY5DBPZx1PlGsaR9u
tMQgfZ4Fz8lwm1SSBXAOYul2TGLkJVPncq0E536MomCKFM37t2KOn/1mUH+XdAR4
DwlNwdpObQOtTfqyDNMNworXQRCd7C6P+ba4qhM0KmOJgf73GUCU3so7PYFz8E8Z
hVOyTGsKKAb0nE+DH/WBwdlbXGI9xNhMhtpcGlQHwElP/cOvGb2zcxKQ7RxNwm14
/E6lM3+EDcGAWUXgR2XktqaheTDNHszjuQHbBOVw7yA0+XlTTv0aQ1c52gcTGIuQ
CupqF1jHdkjmg/3hLJrjtqIXHzBHh1HuMaP/hJxkiU+NqSQlqgyFFsPFMH1LbuNr
w//L9ewMDIW+8ueewB0XeLDV7IyDHuf70a2FSHSBuz+XikArC9MNWQliH9qdSkrk
qo57fxAqFdT37SVYNVvZ2Gx+iCi0IrxXVAcyx3My4/+EeUbNP6sDuavZfO/6ZsIV
fnt62yXUmzLas1atTyscingVEOsKveQfw5NqLsO1l8yDNoLgSD1rmvVIviDBhidl
VM37qNs5AYUEas9PMJeMG4dwp8zJfq065XUdCjCqKz9OX8S2X5UfvDR5SolHwW34
VkmWwsDkuFJHHs2N/40HwWYoxpbSnvEFGF/y2DXc38Kb8D6mU/r17wcSPFZ2sj6I
MHQ+oo2dFcK6Y8lTIBelDthdjGrV4VRPmc4hUizdcaaxSJoPXJCJJ16W/5p91B+K
lCm2buQvskIISX23bgkAgywug4G9TBdqs9DY/YixDjYbNWXmVdj/cvIvOa8vMIvl
wQ22CAUmdXck4Mz9LaA038Aa/cEphYLmIq4OCioB3lluKlen7K74rX19T6JbFrD7
4UMr/8BFsHoV81QQyv0b6HRS0sex3E1fx5RB5fXWHR9fyUX6g+QQ0G0XEdSm8Ty3
EUJoaa/dL87NBJbg0luIfMPHuu7Sx5HTRvbf2s1ZVVLiAbotYtr1nllV42wH8/Yf
xZrn7UqSpLf3KGKcKtZC4r6cWmArHdh8QnRKJ/c4h8TKgxpd7OhJwkwwOzd4sYY6
tuC6FhdWE29hLw2fg+ju31ybFVC8i4c8X1iD5JgscULBuBN91/+ZYFJSNaprH89o
oMU0a5e/+7OfEVDzA3FmcbTnakwwc0sXYcgmbXJxqHDXM6m8SH8F1hEpwC8Lq5TX
jRiiapnMTW3iHuGrUv4lZ5KsjBiBGaqFuBTpgjsx2wRefC3EfPSOU3Mydax1uX0q
HUyrNY/c7sGxWoT+IbrL9TgqWuMLcL4CHemTwpyVycYFgr9ukW5bBuRj9xfNvDnr
5RW3YDhhS0vBabNajlQ9exs6z8bRrZp5UlCuejdgv8beGhRboJciLEElEKE88Ek1
tzMvcLjmgvycnsBPaNpT4JgrrwfJiuH+x6LT5q0YSZCyNMW/lrWHGsi1AP7gXybF
aut1K6GEH9tyLHu3xa4rqpzQBthNs4VlSIh0/9s6aKBKH7NscEfGFGtfjxyFTaKX
G0ZyrEGVzBRwUCkGFf6XpZVetG2QK12qHjf21THahoVVsLuhHmkQJ1EhyNhWiBaX
2wpEa7bhShVY77qxsgCVXK0KhKZ+/aQEdIfrQO1OToIsM/gfvDC6/uM+LEoIJt+o
n80UN/5Zdhj8GneFHoMhOXA5HXTM8RPYXI3i9+xYmy/VTy9StEM+2IM2y/lfiMxN
MKTup3iQjsj0xuIzEHpvD8AGGsCFd9aUumJ9D0nlCcrp9iIB6nThUpFTklt2qkav
Nem8MD6h/I8LAqmsuoblwbur+mUcgUgGnuWKG5LmEG4rRoJ3t5lC7rrgUJ1EtT9Z
yXFmxVCf4PXXWLlpqU7OIZTKmndp3BRqiO+WYM0LxjTRFg4b6o51AIUWP38iMfCB
Mumre95Ab+gi75VE+/uHQ4QQYxlAmXAUGOFY3yDYMf2zrcZKpBx4Pr97fEIjCiNP
g8gaGZ7d/8qkoX/PdDnGjzQAPjgbiRM+TpjGjOVk8GFe6KNUYA5oXJPqjCV7Ci+f
GOXnJMpEItZKPsvg5JMugmyuDJqvdTNk8MSCFeWsanqAfEfXico5JnfMprJz7x8a
poytLHc/gAgw5Q3GE9Y15a1fRen3SmCXGn9NE2zBtXFjaE5RjW8z1aDaCPecs+Vw
7EvovRA7QOlPr+bGRU8IgY/2r81YfmQD50LaEn8sYRScFut4vC2lKK837BmzLrWj
OhERQ2wtyJkCgZJcC/XYgOttHXyTITnPqh2g3ekTzNqs1AQBsf38LoaXmQah5onH
WxprXmWP/E5Q6RO0Ilb2Bgdsw1I9I1CS91X2py0NPSGQi3C9oM5S/uswEO3wQnCr
d3RMhMtsA0rFkW553D9X2ocCVwzq3B92ksNx4hUNZZS0+o0a2pM6vLn6V6u2LVPp
WsELMpqdvAfvePWN+4dohh2DZdxYEQrbprrNca5WZviV6q59meyAnNkw6qZ32IPC
f50sZwGFX62bhTCRpTz42b5wdak57c1TRrjHu2u+MgfXHljNQ0dKJEVMjd13v8Ns
p2sAQGYkf0oG6e5xEVSr1sGwkxBJpi3yZcLkfVTrPDYilw68fSVS+1tMpB5ZfW9c
9DQnsGlyK/IgHGVaNXTs+Ick1ar6FapIe0t1HMIMwMwc8IqaQhE2JPJJxaR1nAa0
Boeed04A/oZiU48cTf+LJqZjnOhtEQsYGXrqfdfke+V5qX7dLPZ/8/CblgLnqlkd
Bbg4iCVoAZzZxTIWQPH/9R82rpjJx9t1RMle83oyCbc9hPpfrdRzo8SY6DH2b0Ga
EM93AcnFitH06in1UJ0dmc5BYSgIYQXu4arWjeLpVunOznLhx5arKq6yB7yLXUOo
9K0QFbhgV38w8Q29nSoBt7/ZHNvlZoY7yDeGI/5t5fXCoU9pnAqKGGVPgU6W4BNs
YzjsHPByjfDFFlPC1owPQEYExSZxEm0KoNU+LuLYFIcESJiWLhSFMv7GKxaDxJ9o
o51tD3HCRuKzOpBpJRxv0i6bERWUbyk40XfXhlbm1B3rMqQckNydCJmRIzHJl/Wi
NsPI6H+GXiAKg37sGG2qvGDFQ3PvEOdGba/YjrKH3AfPYt+7UKqk0X6lf5FV96lf
nKXTUQ+0Soqi4jnmhmyOVvQGhI2up87Z2wjG/mvqfLL1V2jC1EfpjOG/8p9n8nUI
f6O764rUSsivCWLgNLLpuvu94VMC6Im+qRXkr6fjpzyMWg5UX5DQBWxLf1CXtmTp
rrDNSC22AlhcJo5KSa0DE1yA4WjB+1GKLiNL8SVVVvK4aBZhVydaLkPG7Ygy954c
Z4Z9gfs0v9AmbKlQsIylTt/i/cFXiqeq0moK1JEJYFpuXDiw85OkNmVjYyCesBc/
uuwtUfrnA4Qd2EYNPX465tjF8CqGEABpjHkr6BdZGrowidmos5b+6914blKFKmvV
CDigYq0OVFwPfSICu478U+3xSm6mzC2ij1kyX6l7q2LRxiw/F8XYtz/8Xw1PjgJ+
xNGIiTc106h6lZ0Yura9SVwReXOKOTMfKeBHbSWIniqNtyuFefSF2Xi6Lycf2mx4
8mAsdm41WjcxuN6SEm565CkwY8kP/QNGOPapjJcdPqLFdyt1CS6voFBQzACP5qgd
U1fml6caNwbnY+B2LkwQhQjgtnOGkwWbblstlBRAw9cFWuHYRFTMmLDWOoyilg0J
5KTJijraoZYfRCqAw55NPvLDfxZ6HSYPNMLx6mOb76+0VIuOP130HvNDzcIArgTp
F61doeaCnP2PDDXGYc1LLJ4LLT94nXlIAUusWK8D2DC3atfWYaEb1uiUtGQF+hXe
G8bMF1L5bm0jYuaSdQeLMdGu8Qb5fUE29wEwb4d3/AWq88AlFrXmZJDySA+ztXGe
dTwhdXTGGyyuyTNDu1e4aTgt1NBqzWr0Ue34iKQBk5ybJKWNbbkqDgWPLi9aroHY
zK89I7269boiBq0Kyw9STNCSuUewNE/Q+fmszXvJrmvnQ0zfh2nakU3Wj+m3eTyJ
DRlQnfqSBSxhF7q97Kf+Lvq/DlSMhOM2hCTvBcKRqJYBM3Z6kWHFvV4AjrwJ+vhi
rBL0YzVJ9tulXR3A5rcGx09Rcxv0ZRzTwOVZIYN2pdM2EAg9hLXJOUkxkz+KGHgn
6TGpjJI/7P5Lf4bb++AwAT6+pm1VkOXFh4uoQCZlv1wb/X84Qr3f3T8RXeNh+/oa
q+mlBV8fNT98WpxbotPnbTAnE1wFvj6p6rxSLqG+Esw+tjvUihXo+rx1FcSEz9Y0
D3CU6VSTiZ5iJ+fAs34PW1k3klwjiWcF5GtLn1K8v7dPYuLPfoAl3vipn3+W/BYv
GtFCin89JRYk1KhJ4Co17cM+Qv1aO2/fan4cx622JcBm1wknARgLInm9ccHGLYA0
GNbRqzKCvl2bLYacf9JhCqf05LgWZn/pJ/q6Df0p2rccxJagB5J+KF/4+0YMlCJF
i9BlN5MoXbrKUxVgbAbO8WrHsPYkZoXmyerZGIbzbwH13bAvKvVnDOcnIjzrMIhA
PV+AWuZDnO70AoQTyQwyZBR+PFw49lgE+HHFSLqDwSG/GDzLY9i1djt5ULqj3Lol
tJrwJiquesl+zDV0nzvUW+DBM5bO1LgwF6iyxCnddby0nQ8TCIH7isZLLmOUufAE
Nt71VE95QIgp6/YQk5waB09Ed4JsFDMdtdLwO3Lkmsr5QZ5IC6V7uwRt2y1ulO9D
oe3CoqjByVcaqPUGovoj38StrOqiPEnBAAkGLoo902MFZ3k89JjZHCw5baCTZ2Zd
/4bqTI5gt5IeF83q5c4y3gC6b+yfRZWnObGM52kaN4veiuHoDExye2kYk5FCG63D
kZgbMrXC666haAjjrB1xWBOyQn/28/QMDXEYPNqQWD2bJV6v2YdwFTX0TVj1CEdm
qP+rbiEXJOVEUUjI2mzZkWO/x2OJ3RtSqNKcNe5jmz1iT2BULlCUAchR0Pjm9cs6
2QrQ9osAtBUG+08DWbMZK5Bc401pKySMAxFODcwTUjwUiJTIAqx39D8irpa3oBG0
P04ClnPAg2HO7MzhSbvsxxxRWPOl0Wd8Uudv+SZf1wNOC07X0rpiz1eStQGNRdWO
xuIQ0lbOQv3x4J+a2bwOcMhSma3nqB6suDbVhi6i7Rtwom6FUPvIsR5BenXj/sCU
euTX1RCAt4sp+LuCH8JtCAZYoqeTGvQWLJ2Lp5rba+M260PrQUoQnmgLiG34fNBu
+H++SErV02w5Ydy5QIVS0vnjlzpRsZtLgnV58YcraEuhDL0fpKauK4UwdKYNG1DX
KH8jNLOMcgif49fP9YFJJa5h1Ws/XerCmDOsiV2Mgr0Dv1Z5DDHP+PfceCNzSIiW
g+Tk87K0psqtElOC3Uj3td2brc7c9ICdUWymYuLpwfRfj/4CamVL79PY6zXI+RVz
JlVLJlm9xxP69CFj1uoB8zyrWZB8RQsyOb7rb2UaMyZUswQSLXen5+EOHFY/R4r9
gswao/LE87pu99aYVn4hUEHtqlaMkDO0oIhwciTb1gydE79E9RsNNN7u4UZ3k48Z
Mj19ZYLxHQ1878uAfZvJY1pCYNc9eH7CExDE5tGOfkYHG2ZQWbcizx1G4glAU0jV
8tvnl0MSaVlEi7RBBO/PopU/mVArWPeqbPCE+6Rcxb44NJs3jhJHA8+X7Pw2WYK2
Db/ZJN7q+jw0Vghwo2Ijb0z+x1jtgAtTVQz0KZGmt0t1VWwF5lKC3DpatwX9jWZH
fy0Yiklze8ydeSwJ8rkB8S9a/7pfV4mxwanloYfi8zDUhsnrchueiU/Aplta50q6
9Gu9nzGxMzUv1ZBFrhBe4QNN58vA1VkFcy0D74cTBhqSSgodEP+fXUecn2VXLOyV
eZnui3sm9aA5oCEIT9e7upIP/feC5wdkziqizZ1nFy8uxcVZAHXlpU58wfGjXHX4
U97uBLCDydG+4Fu+NJFI9nVMd5GAdpKxPkmk/C4LRtCYf2SEIZN5VlGjK6xzuSko
QLPBhcNqSprPRg/OHQnJ9vGXk827lRmWO02er6tBm9z2A6/Gey9Qd+g0wMczxKM4
J4jGRShaHwELXitdP8yf0S6+jVtMAs3mluZPEfliE6l3TtD12JW0R7YM7oRnU7LH
qLLLFMatY0+LutnX2Q1zKS/IgZXZQW+YRHUE9fYIK+xSTRKucjO5WXCyEbcq8ezn
nvVSLtb1NosOzds/24HS0gyoa565MjU5P/4Rq+UuvfyPi+W+JsyLXiQYirxeAu3I
i/ysNYJN0CI0SPJSztkCcxcTIV1UeOiz54atLGstbMYOK8+u3rV1IGrTz+kJYIEV
K26b9+cy6v2xwfHM+mVI7pkmwWFYe15TR5lzh7ENJY4EseaJnpV7j04c5BXXBH93
jpXFntEQvXSQDPg0tNrehHgGs5sREhECC8rtzXb+WNit6ZZQ7F+HpeizVLXg31f7
aJSWgFsJ8363dM5njJwtN4LuFsehJD5eSy8fsp32IMJi3U2YBKM/M+AFDuhu4mg8
HMkbTWLTRvaZ+blS+2DzKbgoHzMJ36zSOn2ssX5wU9eTvj/DMQB1MpB8/ZakeBYB
el9uY8Zp+LmRzebvRsOt9+NAf8PzSPeHMG7FjebGhDrb4z7UbJGZLCqSMXhGazaB
b1m1ZtEMkKtTIk+jag6K3AmIFwbKn6X70gvDQNKV4fAYsCLzCpRlFfN7cDeiwkNb
iM/GR1xIkFWaFilQPXMJG/ijpAWpGPBGL00yC7fBqaPgRJ0i2WfkkXAU1GIYkeFi
SH5vslFrM5t7eFw6AyNS61GFOyqsTP52gVP6mlycHRLYLFTZUUVvIQebRcxHhSsf
auskbly6uH0wmWphVUreg9oEG/fmz5k92yzGs2D8b6tKsGbHxHrHWpNCQnWdQnpI
dF2KPm8gGowup8++BdydSOYtDKEqidbcLL2havf8f0tqc+5NdrLidHj2MyQabnfv
L0Qc0w11x8Vapxd6ZQ69WCAAym9R45gYBAunOrxH5prvh1DH6jw2kpPJWGWntZrR
e0ElTOPGufdblQLUy7b7s6NT1vgSYynJhIxzaFWqrmosH5RAnCgPfEuLxkDHR9rD
/6Afwsjwse3wUUize/gD9qcmc0qsnh7yHKKaS91uWb/u5z+3EsTGXXBpkg8bBhWk
wD4BRfgSEsAmWOfHNDoxWLWnv2Cl1P2YUdxAO0T9VJLRl+8oGOTq9ZdL2UX+0dSm
wEGCOMLkJzxemCTT/AAiYsYEy5sITHs5MskqxkP6CuKtihc35jSTRm2Ex3qP3AHF
bjine4N7vKZCNay+5VwO1nr5AXbWQGxjTDVWODZ2XK41EZ7VwM7Ag5TmWQmJjWTZ
UbqMemj3Je3w2hDdQrR6bDIuR6uJCeqEE2yHg61Sd+huIqjBSelx4iKi5byAFYUQ
4RytB9vMrqtdo/jK8Dx9sCId+VFbDv9XvOH227kWIUQ/paeybnHO6eWTrh6Aj5SQ
X+nUYOp0GFL2OW0mdLRP9dZ4+AiwIfJj+5nyl1qhVNLYrD3R4oCSR/vbw1oiUOQV
lL8pF1z4Wwj+eBu0pFeOzCJJUOwSCrOgxeWdJPCrPYko3BtMsFQTlGJ3TKmbh3or
HQBkCmELTMe5njGPhys8DVPvlkuY2v4F3AkCRwJj132s130dOoF8T02/A4ToXsYi
GbupvJD/bujO6Vi3+m7lspN6iyxCZ4B6vWcBIOWA4vJOlX8UHJmJaMmXaZj3Jpr6
Un/s1t2aDP36/fQNnp0NPgiIAN75yg094eDuzIaLMKPt15dDRUbHXfXYBKQJT3oc
E7gcCnMxhLPGHy75mKnovy/8ChQyHF1GwccBtxg8ksy1afEutbaUkAoLsYMt3ot9
IXOrqEahychq9JvB97fByjOS5j6cVUst+yLcwq/Ke/ZqN1n+zXUqbpHBQwAsKELZ
rLIZ8aW0olHbib0en0s9NYC0wYorP8huudxbyWOXLy0zLG/th7H5S+MbXDdLtVBs
vb0hfnv5hZ674DX+Z/5yaSYimnGLq2b8IW9E99tC/4szBLg6PuOtMTAFgyNzsW4Z
ETTtFp1O/ZObBtH06302I29V9kgx9ATPbOVKQu8+f8vKtofqcQVWINO7FM52gwcV
nQp8O3PEBMuUHZoTJY6ufjbaEXg2UuItomZOk9hWICdhPz34CIwhkzZLIAbA++Oo
m6IgK69i4N8pQcNZPU9ZvyrKOUiunIv1R7NdJrYRh9xHY+Zf3i+QrjOYDAfMz/QQ
M4ZafDTO0MPE2Qv6kICeKclDfmPO6bWuLQRoG6VbsGNvv7P3XbFHVNQwaFAhyv+Y
QIyaThyMuJ6S1SbzZZnU02Ci4tXphnEs9VlfoRQmDZP9ezXe49IEPTTsq7Oyd4sp
GYpw7PmtXcE8x6Hh0+ZMPQ3amie7134AZjoTFY1ONYh8ECvWU+ocJ/Upf4DYNj3f
faDFFq3LWcU1/eWxx6VrklTSkB0UXxfIZ5ExaDQLf4iEB3F44odz9lN6/h+WzZ8O
vadKV24UcngVjl7vUU3Tjw/GQIQhPrd84cg/YMUsUm8AH20PBhLAvvc6YZz75uuf
z/NT+MmkMJVboTNpwUrs9AnRMhXyPOOV8/xRs+k1DT6mIhqa2eSm7CspS0Axcerm
WvwikEbtRO6yfGm+khqkFBfi8rL576sLSTF8uBlESsAdZ7/rRFGKG2lu+tRlHWMN
coWaJ8Yj56YVioc4mAMAXYmmk+PUcFkcA/yBZfXOHanQXEQt/m/Eg3zOzDc0QE1g
EYY7LG/lT64cKRGzxniN1mz+0nZ35VvzUF4SC9El97Evq1SWVDxsCUTmcLC7unpa
YJ92mx5naNlGIuHzXSpMOFfLsdV0WyFB1QRLPgJpgQMfx2ggLyEp4u8CdI7KJpzC
IZcEVPM1YcBv/idOxI8qk+fkufcpIO2lgMh8XNKcz/UXBVZ00yFzMYsdkVBmom6N
37CWdT6nbgCRc8RVie91IzbUOCp0YegQl0q4G0wLZRgxOwLSDFPQFrlr1FIMjNp4
b6N/X7SogKoF6IWA8cswuY9VaPaUrLXrdzbG4wYnEnrrQelZhRtQCxfJuyIn2TKM
mCfbMvNcHDgos7AylMQAk5I346+RVkvhRBGkzCFWNjQYYEVaXlSIyAzA7cdeboCI
cdSSS/5TrTIghfknSf01AP4qZdNNsvF5DcDAz2tZ7jmMQaj3C9ADt0BAlx9Zv6Zr
rJTw7wHh1I2WXVEa234vamqL7ANJZ4D17W3S+dqNxOnP24LKtqJKOgtqjgEAEvaO
ZHDsm5lytaYANb73ZcG/u4MASkCsjWNlhB+j/NGZHueGklD9FCo40lLotgylK/KU
XNQV4mLzXlERRrhL6+PvSGThJXKlrxNI2TdP/VnUTpQvrEumA+3Y6V/tA6hqcMLR
RUjhh2+GjQWe3c6yMV8fGOzA02Sa0/WwfGRv7eKtE6eEf/fruTyy8+wHmOfFu7vj
WptO+BrT1Og56uIBDWgWhBvI7FJ8qiFG16LBsIG7vmj0C1RDXcPTc7iKlLpcgf3P
eOR8Ce8f0tea248gbwQbZCUwYQt9vp10+D5Vjsjo+IzANJ9qgRgHRigqEjLeWGGl
Bd1pk45WN3PGc7qunaiiMX1mQK7W/cl9DbQ2C6QRTnbrqhwMgLDqaxm3Bi/esNze
hAq9Ex9fIgNTvJDP0/kRwcEPhRlDALpHUaYhAMORnokFym9D4eiugnW8V0RxS2OV
hoFD58U9cgf8XmYwg/SoCYQHtdbFX5TQFz2MkhTpdBs463ilrxHvcS5Q31/pF0sL
wHIRY03Iv+IkDq/9tRIbN+oovTJJKi3Yadqbt0zNcz/9+H8JF2gGDiGLjiaRMWGu
TY+oKEw86Yl7RQwXdlh4Nn7xr8GuBD5MsDE26LIAZpmuItaIcqm7slUqaM0ok92y
DnApuAD299gkDLD+qhUp2z2snpJ3gra2LU69plWT0Vg4YsjuAhvntX8SFmH0onuQ
IrNwhhYAbpnKdcPe6RipJdiZgzHTWhQjjdb6GnbSVX5JQYCtt6dpUGHW0yLqIQPS
SGaAywqCGqJaOyEIZkvstL0jCiEjwjDH/f5vkwVTfDc5BeuQMseprFYxaQE9NXqF
4qNF8Q+3QC1cSQcSq4fGYa7RQPXwKvIonr8gJWkE9IlEveifP8eQR5GnXSFbUie5
ozOz2uKYSQ2q92aPPCf5RSO/epOJXJbcoV5u+/mxLhwwMpFXP3ki3RlnmJQulLvA
4mLlZS8wd7GhZcPtfczNew2gZTVz/ik+oyoWNnLm8XF0nB5OozV3YpRMTxfYoRFA
+jg8JJfX3/mLMIKZ2pvhW7fIykaz0JX5SPhpD09H+nCBG+9V3nCODO2xVfWkpH15
5Q3TvIGa2YoAIhj1+KvNVuVRoX/I6N2ifCjaqJTMM22348U5sm70JR6lRofj/yi3
GuiI3lSCTlUnPUqTuGL+BS3OAgXbUAuhKyvgbDK4vUp19h+7MQ5xrnF9dvWeFkYX
G8dAvSp4Ra0upCMj9t5weJlUKJnJW08AWn+w9ZWt3hR1LDyUPhPjCN19sSu//qqQ
fx/PU+erQOiXY4IHjnRx62oNTHtj3M3frIOVOfXbpV4koJZIGK59aCvdAmoOrjlU
bIITtrkxEstTMfGvvRko3aMVtrdAswBFIm2lbZPO6NkfboJy4PBkXJWmCf+dnw+c
j3PAIgUYX0b7mw/IMTuNHGCZElFH2Q23ZgJ9UR+JE29Grk+afgT2sx1wPYWhvwcR
oX7gfz5HNPdDKIiF62fYkSL37Y23pXlyOydtZV6sWIzrfWEXa4PatoMcZiO7gcoq
mBoH7LCKFynkb42NQaKsRmvGPr0qHD4eGH4Yi7C+53+3NWOBOegM6qQPYL9Ia+kH
HtkSeaZiXeVK6bXK5fKZxeSPfATlmvffYMFE98qkWnvYgoBrJ/DET4BKYrCt3zKx
cPMF8wXI68rgFBLdtwy32p8hozQaA4YwAPemGb5ykgVPyKjRwatDTzQdrtiWpOtv
TbBMWkJ3xZSmf9UAPjYcvHc0fivlV+ef/6mcW/E7e0fYzRWkYppjuYEd2lahP2ym
i5Kpg7RdbufKzLUTKaUYznPsRcz0UDvsgAUPHajG/QOTlvFzlZDV/FaCTfW7IeQK
uRURYNNWD+tKJ+G7RglAqtf5t4GmNh1iTHSuvyYgpQu46zUrSxW/4K0J9qUgWW4t
M1Rpt/zJ6dXeFQLGU7YWDWb+JmEkd4vQUGfJQw3XsCUHUz4AM2V7E7Li7c0iWZkc
mkYZd9LAma+Kv3dxKV363j8tyouqvJrFUbAB6dNoly9ifkg+CtdcSA81Onp2pO3q
w4OZICDec8U4XzjFNHAG6oqi1wpkTjjSY044pX2NoE/7f0mGKJuP3xZBZ50DopK2
bcvvDclX3FCnuRPcDrl1uBCTw26dy6gRQupsrRZiNPbOtCXXccL6gtXDrzMWz1hp
oI7D0GsiGhe4VWSEzdkXnl1bb0xWF5eRHuCW6noYWi7RWZf8uE6z3k5K+PFYFPhw
tGFFvE2NqYnhQwSxXMS6ERfnIRVMhyhFijft3kZmkBE6JdROTqVddLDY7V5nYSqf
YUkbozG4tn1XiB7t9EmpvlhkFs6znjCC2L+nKPX+pHd41lNj344Cr9XgefTZWalh
XQ17PpX8LTWfanPqBtONAkuTo2RNbrF69tAYmuk2pRbr++WVjyDQn/WEClac2OwT
Hb8MOYS9CurxWmIaKJuJt8ayOr3PUahaIVwhUTxQmo0cra0QAIV/fHzw8aq2mUEi
oCrBdLtkn1Rs6Plx88ikpmqcXJSscWSlK8dDs2l/rG800uXFwRIml8PwMDADkbmi
eVjUhoTHiFGjr+tfJ+sdtjM3BGsUvqs+fmtsrBulE+ABowvh/w4ayVSRirWEFlYK
wanXZuvYFYKxa0sjI8S8AJ2w7/f+PACOLzYn1ziDSSVp59bXIxMLiXbuvDEfbN8u
EdxO7PZuoE5AHCg+2XwFfm71pXPL9OaN/w7by3rVJr9PUf/6EqTYAF32b8xyI30/
Wi5HVA2OSW61OH++k0vGIpTW8LxVYY9wUIgxvdQ2A4LlmmTyrSwRzPWCzhhJ9BKi
YQqWESj9oW8qWhUzzwQrL1UsUS4Notr+JdsdiGYAFN0/7dtUcHFzo5kF0W2AXGUy
01XCept7J8QyzMAQlPueSXxo8qGgVwKpUtCR3bUB3/fbCH/WpCZ16COkyssMlL32
yWGMehP+JAH2/bPizfqM2anIMcc7bQGWZfS4AYFd8wGWj9ryorzB90Bi+05PDbee
HSi5haGFFmA3rjitQfm9GI2YAPkhENO7BJ5dI9AmDwnGH4Go9NSDgJgQrYNVHvk4
ghOb29xzGUluRWGZWgcqNWlLkAp9TpeApwH1mrr3xRV1oPFGNbwE9YAoxra53Sat
KRpWYzYgdbvDpCm1EZxAxrtqKUVWKj/9a4q27dipO8+OY/sy4Ie74lDyUpCnNPq0
2i3jLpUFXvCgf2VcTMCifxu9K54H23Kyy+yi4UOVAXROFw3F9GUs6N2nvBoF70qJ
HVSaRClhCcADpLT0txIBpZlVGKleNhTVrbkwvGbCFQ7qfowNeTrIAIg7K73m56pp
5P5C7FWlvpTbBSrCNGEaGwLDyoQ24ZejZquxV9dVwa2ZErOkHwW7BSnz9uThrBSo
FuGL78xezj91Wr8Cs2E29eR4uW1ktC4dGwHaj5epNYK/BuTCmGFjA3cyFBaWj/Xw
Pn+GGvn1NDzS9TM+uHjYY0PxB78X3KGmhQlHFK7V++ak7sSuNXsi+AfISosRMcDl
wFB7rSUcKt8vgwcT9hruyUX+glhMpTGWR0fYbkMm7aoo/XPT44Slz3vigV9cGNK0
k47gADd7wTZO8mQWmYo7z2X4TX4K9G1k2g4tMGjJeqBCCN86xriarOIToQIo0jru
Wf499RAwomkCi+GVL21zbHU3qRgIyL+73d/F9XwB8SW778L8gCHHZzYjACac3kJ1
8ImOAy9q6vFtizFY6qgX15Uyooi2m9EqU/SF86DTAfkirqzZAXdRzDhIO2UPaMUs
QcivItLqHmJJOlt9MD29bJ7Ym+YsXia+zhBTuTYh4pAiWE9OTA+zhgRj+1oGMazs
bv+X9SByCVezkerU0TGfkdaADCCGCJySlwpYjM3QsJVZ/qYp0098eFQ4ZHWCN3Mm
K74PKDBr9ZseYY5SuWD6TlpYNLEox0WAdhSlNrEkVZEeiFXXempvkRYfZC9J8ivc
WX4jB2aAMGX+yEnbKU05hXg1jU5lkPCmXQgGWeDVBoFbH9eAX3l2jS1F1T8vwh97
7G3PkjKMZKiE9rQyWJHqVp5smc0kMzNKXc/n98S6QrZLEvgLUb1F5x9wmG46M1CT
SyTSIOJLBYTY/7tzXE/EJxMzJylKDVWdLqUZVenR6rz4Lg0feHC7yUtuQlSUZfbz
yP4X83ppW8pfO507GKO6Eob2osJnvZDWL+7ZW09OO4iomJeHgR2tw3LcLlh49cPE
oZog06jzPJUzLlKaue16QaTyZK7a+Byy5nOK7Ed635tbunga1wD5V7R7LeUSdgyb
HN78TCmniinQFEuo4bYRqSnFvIaKtzh+3TIBkzPuX9g5do6uUc8WbA8T0DCgoFx3
gRpOf+cRh0+isnZ6B8ybUksum2IpSijLBgSo5ln0BvYBZf1zTOGPQPhYIe02wDhU
lYe65Qm0xCp2dbnYCWlpZDxBy2V8ffylkohcgiweL6skMOTrdXBmRjihxOEfeYxR
vn+ZGX+nLh75H2StN7YQ0qumQUPm9cn39PiFdWQPYIXRiVh087Mxbam9U66gUlDD
ity5VK6U6wivv5fj2GPg1KdyG3EOHyl3Z+EeLICYfS+ZpAZcI6UzsfdNRYsz23wS
Bq5+P4U+ythfjoYWtaZtUm2r6cA2r7aoiW+qmJOaP0+P5I+cqmbkc+u/5zl+MFMg
E1qES07+DxVM1SQ1fX+SSBMsPCf2aGJwgisZ8HLniKWW4FQ2YZ9WPda/Jikzkqe2
zfIyJs3qDex7/JSoyRe+69fXEjoBv7WElBy6CFvWlcT6WoZv26er5cuY/RNNUGkQ
9tcC23yth6ta8Lo+Zx8S/FJ+sX6TjlAkco6nQBWWH5X00JeFBMrCMrqM7HoWVJQA
7Mb89yknAbV2VzlS9tkAL6my5P8nqLFWyMxpZxJn0Du0RX1ICK1asJ+SbZx+AoZu
wFEzhEWt8DJUCJLB0N8htRlSilXKr8XGvEj6p54awcTGO0d6o4on0H6OhhiH5CV5
G9M+xPCqoc0exkLT8IJXc2yE1d1SXq1aPHIwTGCWrDmdvf5ic3QFDGc6GOIWJtwf
GOoTFNgrWyD/wn5VqoV5ecPfKOcUAAQOoZ1g3yJNSPe4PFWdwsTXCWJJgw5fzjiM
obIyXpG3+7EOy5UrTpVdHua4g/xUpYB2WR+q26fdgftz7kKj7d9gaocoL0Wg74db
QNWtyjOsoUE3ShLWHC9wnYXK0hbGbk/pRYKfVGtQhmgX2Mlc1w2airAKFGxmiYCh
KMnwlWriowrgT548KfGNGDVG7eHITU48GZwo6OXkoYDFZhDLb7+LJwKC412EWGnt
qZezcueggxQv+kk47fVs2RpuQjfBDBicBhe5lS+mnanivuKsnXRKygx5PikjMz5v
qj6BCdavDMTNFCLa+iFjAsveMtb3XIKKFD6WCddO6+qK871nx2CHXvDjbOIc41Ny
9c7P7EYHXf5gk1eOCyVcbF7OslpRYMqsshTTqj+U6pfg7W6eQjwaGkXhJL65Z/QA
aqHU5hxodna7E7Eh9Td6yk+I4hAbo6hE7qVTm4wdnHCxFSpbgzDqYT+a8W9pbcIQ
d028LbbCovMj7+K64M9ptqDbsdyBTP6jH6zcxhuh+66ZBnmLj1xrXoaOW0FRm8eP
KpJehrMKJv4KP/dsHEvlmlyPkwOoeaFiDfgi7IY97J3WrFHVOp7WAMSNiVIK1EK9
l5NQE9UEhUUvVIVQZ4g3+q8j3n143teS2Ih9YTpd4RXymEj+TpkvDIMZ3MgVs+VC
PCIghZiv3Yx3sMhbBfLAkWNTwQDzOTcENHbiQFNalN6PF0QIBQcSEnf5/JXsPWSy
CIpamZ+fLF7ZIgw8HTf5ADOE9qklBDymNmEdFhRaeZnEOqw7p04cO/cIc4v9NA+q
ZAjvibJktDBFLBRUYRMwMGMvN9i8GtAUmwZyyUOTTzq71DzLsIyZZ/gWAigfU6KB
XZOSPYydcjaREnGiF6K8IujgjtsazmSVHjCnfjtyOZn563uC4btvAMnA97ZLI0ov
yrCUkao0OoyR7dEYxOjboFBjHIe6GDHCxlHElp3lK+x8HsKGXPG2VV9jP2XwkQGP
Wi8ZTYhnBgk5qmrIzgvf6uDRAwkcJwALtJupwlmixUfOCwdRYZ4WOZ9v7h1MpQcu
3Wp9xYCcds9AoXRlCG/o7ABd5KBk0vU946NBR/p8YocFIE+gs9dB2ME/kcgoL7Ge
5QzNpUl0ExojipJG9s3Loufvjp290eszHLiEfubJNqOHVZbdB0be6N/7QEG/dmJ/
Aey1swXETbA+AJMaZ0AzmIZ/fNe7++mUmqgyf4I+E9b7NjhwnPsci55m5wtWi9np
T6XSPuqXjDKYR28IgU2RJBjSv+KNLY1VivkROFvP6RFsNDSFPFkF3+XN5ZP2LXPb
BLKZ5o0XEWHX1/fcTwrU3X8khZpJoT4+P4GVyBKs8RzRb0sLa67GIwB2kA4Sn8Y/
TUppLBMpOXmn7uAYB0oKlGVjpGKDdT7o9XOwpP5nFIoH7syvHjfW353GRNhLQ7uD
Pltxxv2FI78k1wxdlkbCGO4hNh9525fOIVrRz7rB/GamhC4PV6tb5BZxAoSqj3Sq
WUiIvI8lsxoIWO8O3SQEq8zV5sRe1f3ilF/1PrEwWWNpIJb5nPU7zwzokQ5IORGs
Ag4RaCHIsPcuqAu7uTw7WnYQ6Z3luD8wQy1+eO4sOFKJrh/Pku08MnBxirGsWVeg
JYONoaiCimMAVZJSBA1cVULLXVBuYpX++dgCELXoEyrHSofWcTjxaE86OLT7o/qo
iYBl8S2DAi9EQmpy1mdrBtbYqGlqVFvdiv+NSez5s715XxbPV/BNx9TRg5WK+q8F
l8vr60n9rpwGgWVZKCA6sXTI02mtV0wu9r2nJPkYwwXo/540c6RDuAJC/kUK+87A
qa3j5qKSZMH5I1b53Tp0IKf/pn9lwz41lzZJVhCPZsU85tdQbk2rrl//MnIYzhZ+
bfeN4ueNFWHZ5Wo9pWp3iymGcKermoOzDpOZFHKfMf8dBLTjsQ5x2HE4NkPlNlj3
Mh4wssVVSw7Bh9/OefBik2TVrRpiVbIEBDr/2Cigw8CyGxQRefuXlD6dFN6xaSZh
ZOgZe3qqlGXcOgIwiFt3XnX27pHwa8RbGOw7NTGZqpka+a529Nt8GZpIO7d0iZ4p
PXBLkK4Re1ccV3YKYf+EiC0LgfwHpokVSgmBMLJMkoB2Wx5p9WqziVbCbAULGNx7
/KUaLp5kuKkBDJS4B4EpKAXMeQEFGFT0XNlCMqxoAtyhY8Yhr6+GwA92cD6vaTIh
+1OxmyZm5Uv/WbLe0KRgLHWH8QBt/xKuwvn52sTl1JBbKnEhbs4LlN3y1wB8xIAw
ZaF4wpKR/ZbWBaG7wO6qhPhjWHLMnEPOE3SjP69WN4hKFq1xZhrUisV9J+ajBHmm
OvSnG/zxb1iRiJ3CZxD855b7JAhXVZ/6zky+1QsRrIORJyauuW3kNZ2j55m7FUB5
BKWNosEAEq8/sifo8ZMovjZr88YLMNI9IDC2jlvSssr7NEfM9yd4fJ+pkvB7QfXn
Ez0ZfiTeBJfomwoju8ZE1b+nubFB9Id/JfMaJBWs+pPOfACbzSSdwWtkh0ST4j6Z
j2X2/0ONRsnfM9xIOjjtWK51PjBU/YJUwThXTuabv+BfXVblUINugq52uiuiv+JC
LRL7ADhuQZmNqN2Tna8TP2ELaL12Ho75NGxCN6z7AQtxMdcdfqh7fokQEAIJL3gO
XMtdnq/isFmeRIYbrHOwLjmeeC0vjKhcHf1afANNqu8SGK1rVX4b5WHcoCSqZms1
nsmsIwO8bUgmoIX5bDgh4S1rHInJzdXAaiAFQAcPtb3ZwfeMrTuv+UgcriJ/2T4D
10L3cXpc/xBkXbri0zGcS+Z7gHId5Jje3Ut7/LhEQspHZsX+khi9Mdk4PKBf0wuG
JupxnZv32DM9lUjVNAkVDDA3OZ222IvwYoN87sEvryDIQpg0EuL/Hw0u151tHNrB
ZdJe4muewj7WxJtRaugfC50kmQB/5vkezvl8PKrcgdfQXlgF3bzafOW65lqQgrTR
VX1u+Y0Z9l12EtNU8zUdDQYWsDcDI8oUEHWxOV3szJ6oilROOKlhGyWYexOd4mth
HBPVTkXNYnVWDLwhimj+lxzNq+meBYaxuytz+kTvLeanGuE1DOqSoVEV8Sn2OfVA
2VOOcUKOqvzOiIonTlN6Uxothhwmt3KU8JA3X6x1Uh3hgi8jaky4xX3NLjf9kcLD
B7SmB9oNwz2Znte9zhtJPlgdKiWP2ARwaqRZzc7TAOHdL4+fkSLjQ7ob4GiHqM28
F8dKg2igmKpC7gj6lzvZdq7OXBFMxpMAw0VqYVtb4pbQyUrQZrkfB2kPfb9bkMga
77vjX30xRvwVcqZTJaufH0097QSOa2LrmyJMY520aEfvOpzkB4xUOu+Pu3vymkHt
wZSmHuE5mqJryxTKOr0CX45PjHzj2RyKxY8ZhvqS4ZsXo+Nn5ZzUzNCuxGeML8OK
sn2S98PPhHr6rFE0vIU3gKUDV4R0PqnoAY8Czq+OBLfMLtlf6qJggHjhaiGqXqQQ
Heo+lp6P/UnDrc0y4NWBDlpcBXtA6dIM8AMjCJxTUpqYKahoa9vwi9NK+YQIiXsf
e6At7iRFS0ZJ4ElwX5zxfKq7KP90MnmqgBB5Yq8AJ/RMyZ8481WBgKqdJ6mdGbDN
EAj8Hx+0WCrIcCJmV3iziJd9VN3fmdfGqJ2nkCjeiYAAEDz4raZU1XP+/Dj820eO
GVvpFEwhZNr2MmZttRYPp2/A37TirTbMXYtXpVPmBZhXJy21w9KkhAnax/gM58wC
nJ0NRhP3mk4SuPPaNGkFADC0TVBuAN8+9OWU8ZN5f6kaKNPXAGQUJMZKHbeUB2aH
yxz0ealRduVmEzfGwvST6QxBZ1QHTq8otMhnough5ZylPkgH61Aeox5Q2a/StF4G
3JGRDBOYucBSEhNGLf7RKaKtASzsqgacQTZbV+uBDLfNbHU+4Bpk7CmDhm+SKYXr
IUot8493NBvbl6bqERHBGf4MkktP5ruEFp4h4g+LVVZNZK49ZIseZQub22nxzpzH
FcQdwT8mPm/7tyhuGsuZixGrU7GEa2B0bAMYVUzoGaMGHuAIpnDu9144Vd+VcH1c
3TqMa3Py6jXpTrF/v/7xwE5TYNKzl7ntndXgLKlAmwjPmdviZQDA0/7eRx/IJayo
mZoRMvpCn2LdCSGJpZAtZ9gEbAgrn8DplBtT9uXfMD8HAmLCBRwyhDAWWyCVE+8/
1c2bYOoxUA/6VWKO8oPzrlOnenttZJMMKG7V1lhIaen5ApDCUl1GlkVCuxVVS4g5
pdMom5gaGsJ4uDbCjrqdcFolj0g3suOZ0vZKk8kNXeJuUlwd5Rfunc2Xyc1P4f7o
L8WsHGiy3NwL2Dzxx3ZfqNCSlSNLbIcHdRt0IQhdrFriEBVX172bJDukdN8u328W
CYOeKjFGvqmH/MdL8Pwz/VG4/Cndvl1/HnpRHyWIgGpmCucv2yVIYj7pweciu4WU
3ouFUbs0Ff/w0EUeXIbvav+eT/+cYd7VdhPC1K8vdHyMcaxU8PdesApIZOdr9f7m
MJ0HL6Df9gVt54isMalE27VRjiS884aQ/FoxNgO0NL+utgsULCHnlEN0XBsHg3P2
CzPovFx/AAYidCTqs3Uctuex2njhRkLCWUt6Mr7yBYENMuiPYQBsKuK0g7Gzhn2A
Tkzp9sqLIBxCbHHeMPxSOGlIr/lFVKPqeKAuQ35jjGaBKix0LUwkZlsBsS2y15U3
isDgB3QvO28x33L6i3x5SWYFDkfgRg00PRZTBpOvYOXWtyMjQxy+7vbJHqmy7GQx
q3fvErQbSNdU3dvrEHFGoqzFT3JeHN1qampI00Bl7JBRnEOfat1+pod83UMhlVvX
DruZVnw3v+9oocZWIoTiXUxButXQTDZG60vBnc4HkTwt+3QzM5yWEwmYrDCLK/d1
tROlFThQXQMi+vY6CENU8UHcwHjwR00Gai7PcBu+faQ3IojfBBZMWf51G7KKtZh6
G0dOrLNFvHJ3ZUgKGbXp7Z6D8kaGCmDNsddPZPl7CbwXLUmvEd1IYtMIIh/jQEnM
S9pHtV8RywprHBgprj6ASExjlD3aTulr9khqsWM9vDft2sMH6HSV9Jw8/sTPRC9I
dG9pPRwWBJ8O044XEG6/dR5cdU2Q9VvkKX8UI04qAdZ1e5PzglBCMNZDN4b3mfwp
EthMQp5SwdIZMLw8xhkmivFUNKg2UQUvXgnks1xcYHHWM7pvOhiU9AubrWVWXLvb
4QyXq17HOdkdXhyL5Otq6WGnsjqD7a3/PnQLX8XBsKu6rUq99Dz/FRxhfqGC77+B
6M6cSIsJk4km515DnPrTbEFVNZ69NZ7nYdwos3Js0uZRGGEjgNELqgwvh0dFs96z
gS3qzxTQc9ZZcOapjuNvUDI0NAPlhPZy28exhYzmO/Glw70Ts88WTFAJorDa3fiU
XUEEPLemVjeO2r9drVVYooH7gnpcpnP7cca5lk9Zt5VeZpBE9UR5EpElnd7mCETe
4s3Vhb9YEdAbLmSqWjqL2ZARrq26CB5U8z6opZC5MUa5Z8oNFsgUQSKtNU+kqicj
AUZSMIuP0FQhIviyEvQyaBj5/8Rp9+kly+aAR5883b/qOgEfj8Yko0Tz2BpZTxNb
nqpirz6zeICi06BIz5YF65iYN92JJk412meEr/qtHVKc7YpWxp0o8QTg7377XURn
8aMM601VgpndDaTT3k/sQpgKwAP0e864I7R2Ehao3b+/yk4pdW6QAL9RC6CwPWlB
li8wCYP0XnRthgAwigx98UIH368ehImgSTiw2J1Dh/ttR3qVNAu4tL5PAcwOC4UJ
qtF0/o1aOBCBE2BCNmbyQxg3Ann4f9jJ7JlHGGc2aMbd+V+bnHrXX7uJUTt4xtPv
U8ffk5haPMxR4HSuRXx7Tt9/3SwtP76EQqfd3JCH6ZW4j3fgTBRP9fHDUWQxXPYJ
TdRRTL7igpzc/gv+deGhWC0padg+4Ewz3MGE4ySQYy6IQ+2L1zBAodYcLHVoo75t
RiivAzlmp+ISeB6dgTgjlnCGabIpDo/4oC9UYYmdC0FXsAnPvG+LY/22TibNHKqT
6vhSmiUaL2HOF2pph7dJtXouHt8JFLJBK4Rgh1K0U1omkK5MMqxQT8dw1NsDs11X
gGsbpbDWTY4Zl1h0KM3SWIWzPKra8aY4yflvQGVC/GJ8cY2JKmsXa4DaqjdHXjtT
f5hIw6ufsgH5w8LlkSOpGt/E013LeXYqNCUeiZzIDLz+pRwayyzw5MBPWYGEA/tu
Xa4lhPvXZHdHlJFC+7nhxNVl3v7IzZJnVRNUMSSUt1sbQoeCHTa0WF5J2X7mK2/9
lYqHTqhsqY8zhokv9NfKy1NZoNHj9iEeKZsZKPXUeWL0slnVg0R+fCakmpknb2bi
G6dqxo8K0+GPlvzFP3Etijrv1t1gMgkdByeXVid59PFR5M0seiwX8VvjLqF/Qn8m
1lLVNGV0S9N6Xb7CGk92aKk8l9KJzKrA8dLRbQWSViEw0Gk0iWdbF8JaJO9B5vkH
SrNjoZbq0Q442t5C6g0EOZHnhgXvBrDSO1cJg6RfMeBEqqqqhcgf2UTVvcHl1vlr
4HQZXPStRab2OOedx1MDCzx6eyDjj87+SqBNdr4Si9dB1+W7EeS6WQlEh5ffymGR
PF66DUmlHMPGeO04RddUiLfx2E5+M2FF1rZNcc4Rr2Tlclv60rO2s7pMYFHsZFg/
yvmwxaDsXF1Xjz5CK4le8ewv6p2kzHCFmpJWKdo18Y/uWjS2n5wUluw1dDdrghRu
SMoLWOeXL4KstY44cNnWWmsDkhSgu+8WM1s/eae+ZBKUrUoj4S36OoMZvtv+tr7E
FeCEMUQfqPN9B+QeZcg4TDRNUf9s80pJ7S7802lpdVfC2rAtMn8n6dra4LvautKS
exfV74kt+QmcJNQZN4/qnBQ5QmkMJhUxeQHmtwmdu+yrvD8d8FUpMzICXsi7nB8r
ZazeQ/rCc74NiD1UzQMERmHiloidrSZgR5G2azeq9vReN+EQyn1zFWy+I1zAHNAB
aGswrFxE6BRXgM+HfQAaXocp7wCgqhuDKMl95aA7+70hnzUdFrd0bry7dio54oxh
iGJPTOA0H04NOM3/O0rZmL9JYX42fTRh2bsp6omItWLJhUeoscZyIdh0j+ORaw2/
hhEN0CpSuRhhy8W08RMGjd5vwuCIhUyRgYHsXT6NkydaJq6r0SFARbDzQq0az2nW
sa4Zih5JyEJ2bHvQUlzWWtlicGcg87JEO6htABJvscC3ggCqZOhxdAeknvQeZtqK
wdeVq+U//Kh7/q/tWyyu9mrwya6hxvIa+HTydO7ka6de6VR0EyllCLsTAH1GtV0/
gMo/mCSIwK6NEsLOfzaTU2JD+KAWMHCnW4iwGUxjbQviKN6BdeSr0CzO2WWiQ+qy
I8vy91GeV8ovIF6DNOz68Hk2ckuGmsUUf3SHFUut9fah3wAErGuLMDk7UYsvlF1Z
+89ktK77N9WPyzwuMSA7rWZ0ZtiUjfukgM0/0YdzjUP71XOK1T0g0xg9AecsPljD
5R2+50JUWgIgNrfOs7b+iTckL/gX67Ng1dNcV38s/6V2Hme5tlxIvsX76K1jO7/A
FqRP0LJCUm9oba5wlQmA8a3i/OrK8RFIbb6GFc0v7Df01QRJQUiYEEwWuFPpLc/l
h3f0NHDkOT8VLtGLNHE1vRMvaTgOFkukzRTv6SG0L65jqcoCZaR6xSvONQvko0Y7
IFclkRWI6+Th+PIdM0Jj200AfVo2Ge5rF78ns5MVBUOBCEq6ClFev1Q/MOe7PA0d
KmeNXsN33ar7RXUEdpoxHAKwiE7919fWR0HB5VrXvYp+tFFAKdVhr90i9ZJRI7CQ
lLEDPyMtp8JPljCuQZr4KgLtJpPe84l7jOUlX9Uff/BXBE2eZ7wSpFTalomG+z4W
5KTkMqaSNFQcUaS5yCQ0uHKkrmtoAM9UTE4tds/U+NBTP1tpTDHCeeXwBynLaeKE
abKQ1xuRokKFKLwehEuyK9kFsL23x6B+3x29f3frV/DkE2NMwJRUZ+NjEz3R69zR
asj2bVJjpNueSCKuroDJ0WbO2eI8hLvPWV/wxMiDYKLNNhAolRmnRYKsW3CXveJh
Ey0E3OXEIzcdyeRei2WVE6QSz+tTyR3j9qaHhWt4DKGsA3LHM+f2MPS6WGbGN28I
thM7o0P8+xNaLMWZGTCZ5aNLpP0Rgt69SC/oE3FHI6QVZlQbhuMUd6eFanbCtqty
TJYpqNkpJLsnCeXKjEvNapKMBWDbCS5sQyExUZNepY1ZhG6FutqIHX+91bJ9WSwN
6GkxKLX8E0MRfzsOTNpao5ngRYWyo2qxTgyIFqUNxiR5Xf1DGCDSKTwzaXQXllOc
JP0X4Ur4uTY8Ny5Yo0hqGafmBFRKLM3C1mrXWKYxw5hU5rNHj4umFRK0pl89ejPL
y2YfncyhJp872zIeZ5YSKge9lUEes2N+KyGCnMjhw13vIW7w/gjVXvxzOBfGYtV1
KaUBvrHyJd5dIKqg4sCpj6wQp9iS/rrJ0DKhjk2wj/M/c7jvAGMz1xD/67mcv2Gi
llu56K1h5Aacslt0SvXGVfn0ktx3i1Nv2eUpZICGxRnKubTBX1pqg4ZUZZfrfli6
+SBv5oWhDCy1RO4KjoK0nfM6N+yPxHX5SKaUlsHTKzD2i29lmHD8PmgyFHdpRjal
n1r6KUhgc85Odav6mWC7majGmb4L0fYgd3JzzgR2WeMmvE2c8m+5IgE9DSiFWiXg
go0ZdEz8o6V4VMFGihYFMrgsNdMjU5FiqJAYCDPRvaaJVOy9Ip7ekDHL9bPoTPB4
me8UYjH+bRt9/ZyYuvuhBa0qfn2jfJlOCheB/Z+BlJ28LyvW63Tw+kiM1AkeF10t
Zlj6yLoz+SO/rD11j4+dMjZeQ+Sr7NmhqSLzUHPvJMpkWydj2OIYBSSicQfjXC0f
8Nv1nBvjkTFA4zMhH61ONkiQL4U2AJ2K7njIl0QN55MtnS+MP9n7iuf7dEv5WiB9
BjyQ9S+KcgotcM519mEKXxDy+ui4PDK+kKsoIT3Q4lnpJ6NoLHCEyTVt38PMqroQ
UKff3arjT1/d7iieNStWlPnE1O+L6Vz9G4+r75G3DX8BN/uq3BSShIMca2rToMMg
yJek9E7Ix+BUZNe9gvPPrdXJLHkVpFUtgcRoEXJzMHKaJWrWpxARSOCHxDLYOURE
Xzq7wdWujjbCyA9iaMYF+o37Ok9k8Gpe2nqWjmNqXal93VTxevzoYIZh5HQpnScA
bwl0cmufNDsJIMAe6D0N1V/BpHMutRyE0HlYwGhspd0mWieMn8widjitJTFde0CL
nIH4lLog58WS4Pxecpo5xTZpAapEZaHJRi4wPiKITbqW73Pv4MgAuEMqpr8M9GOt
pVBBffifuKu7Y2d4sv2ZlGCzwoj2QZPiNpxDuE367gKRooJJxN5iJ1+RjDIUCAHj
pQVHbhMwjDyRwy6PeRawTvVL2DonuwriVo5mtDOsS/NpNeOLlZ7V63/KCXMUKbAG
wFaR+usiK924oHdWDv2GZwhP59ehuLW0CoN0kSuzRAxbcRSIRq/NQINVgwW0RyN8
fgTdtK8ILxSmMypbgevirDE1XOCFW7SSt83NeW19uw2+uDCIiUVgABuXjiSxUevR
/HqnwFtDq/JRxll/wDivvYpcUicUTYKEoNYGHlzhVYNMpMEa6zIULlNE7gpVoXkN
4ve7i0rrKHc/m0mNIwbllj+w2mBycGaWDfS+2EDZeUv/53QmcfOW8zBHHyj2d73B
SPq48iSDTjvHaqIqHWrY/KYtavUMrz7Upp9jSgXgglpvdaZkf16yVakaz7JMUtvX
r7ZlqlVUp3Ot322ACRztChWMiiOnCB+tyVoV4ERjiYf73gBlCOiBSau/dIlwtw9+
cfx48tL6kKu2ifhQmi9BvmZqfhgkOmg/H57fzvafi74ixSuYdpdIcrWsl9eZKWXw
+P56uHBI6+NP3vT4Qk2PEQsFJHMzZUgN1W/wJnRP/G4L0NeRBTvbCUQAYQIJo3AS
D67F5RrVakwVTWfHLgQjKBK1+6EEMtJhDuw0VKuvevcHYKiwCrvEu9rY/Dodhyfc
7Hb/w89K/ONwL7oJkJnl3DVDHwf0KfuBnExQcHNVfkQvbZ2jIo+GWeySTiBx8rQh
SREyQ+QVv0n859b2CuVfWzlGWTjUXdcVXdMxluASes2DmWLb/1vpf0KKFSY8XWKe
03EKlJyje2PEXKa1q/oNOdYy1jMXm1p4RZ7zbHlWmR/gjR9DHQPj4/lFJFufTTLZ
xDHMG8iye6wyYXCMhbYSMDNv/No5AXLt0bF+dvC8hx1jjKyFTutiuVz9F8hpN2my
cd85kWYRk6Z55TIbBAJFt1xK1AwF8KpdIHdbtr/uFVKawaUY01721G3+vOFdp4Gb
AG3JdlkZYapSDTt0wvEUmVvaaHU/Ttw7hUfYLeETdj9NYN6dEjf8Mx6BQg9bVFbZ
QFIk5txKqHsA9HVmP84M7LsjShbjZSzc4RAnRkmy/Jq+Ob34waBueXwvmdgYiHwI
4nXwFE45ElmEY0eU6UPeNDRp+HMU2jq1+7diuoR9WtWlqGAphJ7REL+KKCA5ar93
w1SOP9ZAVJUPOoX+h+ayrLp1/IaLvTcQUtTeEHZu+1r7bnz2dpIdwhwvSb3OdYUx
b15Ec6mAlvAlJMLAvNppfyQzyls1iDcBW3egkT2Ao6S888IpJ9n6C6M3YOK+AtzE
EwrANXlZQgt9lcg2Erk3hS5tuyVx57UEpzG3LxThqDr4HNixvW1TzDSP1WvliQI9
xEinh3ldrNuCgLEieIHtrsZPg7n/fhArfLCbx1xPQfbjjLARUSV5CteIIHOqVSIr
Y5dpAa5q3Y8nsx6+/4G6yOBwqgRNAurhr/W2JPl67RRBPLdorquFx7UiE/p2M318
7Rc0r5/80OnXeBii+ATH8kYZRWBgnurbUfkQE/ORmlnO96qavbjYzKPG94mv/M9A
QRi1OTw+c5lNoEaR0X5L9CikB5IOMRMGIztMHR98SgZbNqHfDw9tc6vXmndbDGBt
KhqP5st/PMMtJJPCAX/0X9M0+67rrJQNCoWRRC6cMnERXm44YUFq76J122rNQpR5
LIuRe2D4Ofhd4oxW45NCuuJedb29x+k86FCSe4WWz50AuAN8/oL7R5FQpIpd/hih
N0iPcXSmwxPdz/pDP6xIkM5qFrDxc5zVDJ8QHtLRZxiEJOuRm0NURhpGpzcuusxs
BFVDxDL1N5Ovx76GSD5M/2lBw8Qkp7IngfHtYnmP69vaZhIxIp+F4LeVC5aQhHff
tearcyFzNxOZZ7oMfH6mv77CxrWe/Htcn2X5yIcK8jVi+6eWxFCmox+MlpFOT7e2
K8MSDi5PPzt3/62jBcFRy6iYm7EDCDr1gf/ZZgNgoilCEuIFruLDuIA0RJ7fv8Bk
dXFMzSfDRkfna9dOnRgEKRQD2IDkDuuSlIEGfBX24sfDNGWWFUUzJgPkRE3Yl/O4
ZoPE2FHVYAX+7FR8NptLJh4ghVWVu0H5PLzteTpKHjSvfXc+8zqZbZey8ZuvTgFH
dDsEQX79DBSzbgSaRCys0b4uwj2Uxi9GYCnRSTLEUucR/SngTb7oJRd616zqQAt9
s+68waRVGQJdlnw4iSzIwPWxSZxrxJV9EYOmR/cQEsirdvxiff0Pgd9g0LSr2eeq
Ybwl66zVZ+0raA3XGn1KwkdSS2f9dJO45ESDEO41vp1wsk9WUnJ7za+cDqQjST2q
zh/7u8sS0gJa4Z4eRqNx5bSkOdt6MuvtM/4sU12ilt7pp3a93JwqeWmH1l1n7agD
24OG7kndF0/mpW55OIMQUklEbb2HgnfyLs2tTvp43O5wK9GnNPYJwz8rwCH4vZ8n
vZMrrfF/RdRet6tqCda1lpQoUzupdSKWKFKGgX4iDTJWIXfpbCE9iP1ANG5Nc28p
hFSYJtdatFiACgIDC0bP7wjfM700zlo0iyaXxHptlT5yhaKNxO7zxkiJW8c06kBe
szCtL1ewXIhZw1WQtdAeV+hXyBq7JdXdLXp9RSxYFke6TDm5OgNFAxUgPuYjuqD4
EXzjKxOyjRsFkcxUj5fKN0YWkRKz6UCxSgshIDX5aj+Qu45x+FG47dVo3cBsC819
VKLq/hiUEPt2VuMNW10UehEhM2wiB89tcjB06t9Ri0Drq9I+nv1RwwcokvtGDe1s
mKA6RUJ6yWbrZci+HYWGBsnkdmMC9STeLzIu8CJu4K58rxjygxRY/xwBKId6SLBp
MJUHF2CWzdUkrJBhSoz1fF0Agsq89RJtPSAGKS8duraARxO9C6g08WAFhzU0wUp9
mlkzravpfTWuHbHYBEXaEiTjS34DrRk28xkwjRR8CZDu4Gz8zZvw8M5R4va2QY+M
xzCIY9ggRd52+HGwicWIgR8dyzj2k4VqXNsomPhex2RIFGh638mXdEf8fs2a22vS
/kfryxZagMseM+LeiRvjlmb9bGqIBBCzEtSYCLg2RD0pnTPJ4/XanpLWTa8KP2Vq
APECGHPLwXMNSAC/F4XMRUSmbZTwkHQTSYutI6LGxD84+OSCiwGFMmHWh3bmBUIX
xQYLf2JTokSmq6I5kmwNo87kwxP3GzIVxWygKgBu00Il/gqMiTEc2vNkVDqjMrIj
LkDz8YmXb/nAbL+vAFb1RPjKCOnqugH0r9zLGeNkgRHXObk1fgorXHULrchB0ZmC
tTQ4CNiHfww/YfYBlRGCYIiTPctBNgHXaoOBC3g39Xk8CXyXS1nt92I9J4kh7PW3
ZF0ZV7vlzVE8nPb+aitpEQ==
`pragma protect end_protected
