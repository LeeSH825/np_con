`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PQfdT3jeq2R+mreHqVWPiMF1QCl+jPxmlDWP8yk4bbE8AzmpfKMIAXYBcUzvF8VE
+Pi5lD33Bye7waAUUlYhF38XfXumeh8UkwCXVe1HDsnbaqY5Vlc/1iblRv5GUkIL
nXm/Ox3mwPgPWyAaotOwVpUmJBseOY/A2uTZsN+YP7Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 66608)
x3/GacXRJbOldkzR4baFGmU/4N2BIdZ0gy7i8Q7BGlM69ZCn3Z+nHsmtSm0N4nSd
Bvp8E88m94aRDKGVUtfJ2KL513JordGpL382H3t0dxLb8KwWeqjlu3jHVS81uOQV
qVF0NNVeoqt4vaswXPMXMZJzUWt6ayuGgUhCP83TaTsEsG5+Yhac19Ddzp1VxZs8
aoUe6hil8+J4GW3ATGZLqQbBLhfBUNtIi+UrI7RnWGzIQRU31qHZ23tZXEwdYnCO
zQWV2JBbgMzGbAvMgWurYmodF7CFmz+0Aqs8967M2Ao8aKcOfeIh7s23bqjky/fR
qOs2B6R9UP5hMB+B/AHhaHPPeRZkFCEqmaV0PhwsIgAkfUjJ2WoQVb8UdNXywasf
Y5SzuobUM3DS1vABdNYv57h2VDf99pnYfKMAUfpmxFvXeA+FmVC2as2zEkr1Qjw4
jMBL2J5yARW5+eIC4ZBIJhgH7eMorSkRK1PoUldvARbOw5lY+FaDafKRqgFWypfu
NBR0JOLzKNkjnzebqgIJ46mz+5pD358E6q706swgNQMXqSKUbekVyS00s7JRlzjJ
kCOqbTr3tQSrlRDt9zl7ZmdNbBI7F5RWzo4idS04LNKLfq2wZwY+fWiW4PHT0hD+
i5ZXANg9pyku1rCBhXSb4P7xr8YTyOImMKvJ/WgljEtGGHBuTHxu6vlUWrNrLz9o
TVlMjrpSfSCxQ/IYywnUXjf7nej7m8P9smsFsluQGzqcyQdTnm5tx8HAizXT6oiN
sDdQM7A+8CxNw0+bkWDh9kSesVbbyX7aPDziZQcgAGgFIfGIKVGpx3Rf3fxdIhCg
F5DcyuOxBtMAT3E6SCxOu1aDYIEJxmwBcyjhiIEajwaauRoAw3jjSONybtLpKvGv
7uPtULvtyOamWiQsEWqQTuZp+Aa+so+DuKbYtUJq6ApllwilkEjpk0eNIAW5I29H
+XGMC8pYyu4Ac1Pl/5P/mflIrdidfTPGZJLDeqfId07Cwypb4qd1h+d15kKoz84d
Tc8WAEXMbvoy9EfpJc9Fd+DqZc1KA9QvMzD+rhzsFzFiW8C0/kfoiPpJZv6VzR5L
QK1OBAlItffOoitYyDPKoU7tgzXP+3sDU3ZTz35slG40hum9STHqgq9yOx5uc5dv
UkLr/eD9kQRweCBsZHS4Pc9z2cAtlpgTevgH4q648NV8cyiyOUDvuLq9qMZoB2rJ
sx5gJ/w5OCGcVnV0BNEmUrldbbA//WI5sXj/u8xYS9BwrRMNFWXuw0eah6+uoACD
Hb9RLLWvLy9gB2HmQ1HECOKkIH/4lYFNtv0XKuqhgoKbu0sUiK0Tue54VURLsyDz
UANlttLVRSNnB7VwBQPpJU3QB4isxJQyuswSAbnppC7WUDp+yN0veBD3tmfVTAC/
dsz0+bdPcwZGtlXUyNRaSQan5R2wG2i0LZnyLBNCAdSK6c5Tfk9g+N4+B0l3rXMC
qIJ6xtz87naBs61gS5WVe+xTG71Qjqu7zStZOd3+IlYwU+05euVUjJfH/mG2kmcf
4BnNpLHU1NKaZb2EY3s8E6yVSYMwNtyd8yxtrD1SKMW0zKpUSG+WQNzkBMnOD0pM
vknaKu+OjOP1JPkimMb6z6/Kwb8b3B/RvhxJ0FCoU5L1S6yyZaXGAcLzVxP36fhh
xDlpZogFcysdf6Imj4giBVFcHFSHIwIUodtxkTmmQFX5boLdDVUZ9Gh93BSMgH9Y
jUCSOGVDANgzjtEjNaPpCHAHG1H/CCMgiC6t6F4tc6Qqw3nbBvzqPRv9CJGH1F6z
XA8sar39U0Y1lk3ztAlHvRE878fc7y4HcKYmHgcQ2EV2eCeq9pVZGTDUC4BYS7Rr
iKyqdJLqC74QGV/Dyp75/i2tFLdM3DmaHSkBnYvdFU7FsQVXEL9xnVVkNwQb21ot
UimtsKXoK7O6bQrlYidLr30jPoy3R4Xi2PJGzuPmIeqriiXnn1NBFuLtvlmxiK9P
BBzquIDBhJ/j7DsAJOq70xI69OvKW/nU7g8TD/NXCVgh85t069Uc6q0P0ArU5Zbj
15Rvv3SU6TTLDxQiFhFmDbtLcMz4Ye21DXmE63mf36RaM+xJJAt50bs6gFadReBh
ukx2MEmVhrgajBi0F9BaNDSwlWGF7UF0GBzCciQNEfkQmL3mocr/OTGK2/kFxeXE
U9BJRf24dIVdDNued+T6gMZCAqtnZSaVwJ75JiG/zY+SpykOQopVezRh+qUnTOOv
9f6fReK+iIA8DVtPeuBrV98CuMK8Pu3ti54XVsHSF+vBMd/gID+rCNanAjjqsf+O
liabw5i6IfoXwfnYvoQ/sXAIPbouzVCr6vtHuRVSR9PWhY/1aLCZPZ5EM4aTkgVx
4k1cATykYsttHzsZeqDv4IFvoaEyYRmgHK/AhDPyZpcNKBvNJkkq6fTSnasMv6N9
inbPO2DTPoc/XlZTbvjX+LZyklTCscN1j08zuoO/SM00xS3m09/sYCevpcX57HqB
y1wOQ4L5ityqtTui4k4AjVnMKuF2osdgjwOWYCJp5kJAbGUhTJjsUFU/Q2tH6gQA
Fjpeo3bdlCwq5g+Mx7C4w3JStXbz7wHwJR6EHvB4VzDrlFLogwOxU4SmlXJ6bkOC
ULzeE8LOQMGK++lys2oARtga6TM3rrVPvAFC3O7xZRYsBs0nl8tLJxqto2OblxwU
JbE/HzRc6yW/zbsLyLItqX0tx9k3Ca4iWTG3Cl7oRPRfHk9gDDKMBjVvLswTDkeA
dm6YC8A268+gHSAiauPKQENX1OHtU3mfFAMSwGwjP2WMELLosZhsXCw2cd+T7ayc
9NvHPv7LETo99GJEFX6KKDxTnTMi75vQw/iyBbY6FRUHSrqkUTmulgk7f9uwWl6K
Kz9nXWJirBT5++wyyg6fAz849Jv77hkMQkjvil4YzomYMxId/fOIpAu5yzlCMCl0
JKzl0Ibmhn9xmYR/Tpn/3S4BdXSzkibm8SK7SGbvtzc0DVjZrFnnWZK0sIoMDEK5
TLrqgGtmgm0EG3uU6W7CNUZkuaESUcXjolIS3oeuRyP3FiaqdRsNF5h2tescfWhp
xVzRaPaT/r/l3BJKJeREKS/6PJ//apB764gEvw67Ir9NeOTqP9OCv/C39yeqOVa+
24ygQMz17ZkMiZ0FeySRPaZounicY9MUra3PoVVppsJY5pR+WtACy7xjFp4UdPw2
ofuWtiB/tbhju4NDG2w9VFaE6p5pxt5pv2MSUlcxzNXozBjyL3u4cuTnNif7le96
L3P5pEZXOgG1Rf1d0BJP3UzuaZP+zOVA9d+Vk1ZFQ3W7BH/EURc/ST5cJj22PIfF
yVABAzp7idg+KQgo2FrXNxPDXQrl6G9o/spnmJHmP9TtmGUT6xWS5o9B2wCG6Bt6
HG56DKIVK1Bst6SEfGySC3nFsNCXQ7AZIn9auh4jraLrm4B7I7m88ivLJLEhEVb1
hyPZyEVnBhd44+bGuyasjAkVaipTkVkVELdeXcZB8gzJ0f6TrlfYTS4YsBN+NzqB
d9l9MoOUVtBLPYLLvKWx8fhpRdc0enTLJjqI6OxoyCrlNcFONPTACDOzADX9YotN
AavWn4WRJKuORCib0yXB9XQfuEKqgdYRtdV/PvicEo9E5NN9yRqeG3yIsiGicY5f
2wP71Ut7VURG469vo/jTiCLLK+9rp58dP+XlhWF1pymExv7Q5t0BcSZPTEmS9WUd
xywgsZlGhaxdFxXwlsbmyvVGPnFAUTzpuwkRRtHD6mAEG4p+bhZWeBl3OsmXFn9j
NrO1mxXRxUBm32Xl96myGXxqmpUgRLo+RX5VG01jGuXe4Wv0DLcNN4P7ulXiGaVM
kWs7UHak3u0Kcnd3Yektit18WbH24xTfOsjs4mUR/yNVfBJG4agmP8tyHMccQ3dU
QV0+zGjX4y2j7SvXRG8K2MA44ei4sa9dh5KuP8GtHfcoGeNOuafYBLyFWQS1Jrbo
yAqUN96mt/s3I/EU6yWZrXyi1k+mWgd1unyBFsPQ1/tUi+1WbJPmPAE7SgajIDtz
Ih/QaAK+y2EMVYmMtdgEinCTLVQeswzzbDhCRP0uSORVaOwateEZiDlv11gk+PHr
7PX3YiK8WniNZxZDd8pcVPG7/niPkBJxlDFludbLuHBBSOxVgTpaUAzTVQcvflUy
6LjrlF5m77gkaxdqGRQPfGmULs0mRLOB+kva7LEiG8desMfKDXKdiWBXNJjI389f
wF8OkYKAG73Md6keB3/1ZFdt2kDdnS3gOd3/N0Xl3SeEm2CycSOax8ZsCEmHmihY
S0ZYtTEc5eTmYvuEySUt6QixTSm/YjPVVS02GwIAX/VxnG0yOYSblZMbxBCPBcWS
s6HuE2kQ6ItPFyu8NUnluXq+M3lYHkIh7goFDlfXQLCPR0Jw5FKLugwfV6LLCn4D
CGTrOIo+/kNM5DL1WwmSxiFBgFA8W2M28Vq4Wv2wGPYSSbSCYEMxYPKhaIVtHBg8
J0oHMR74vp1+EuIQDKaVBiVRdS+dBTzTS4OL5vJwWdDmrTp3SalcDb+U2a0DuYVX
NNp1UcRv0yJu6WYGg0kZMCwVzoGoAS5FIbL1W/idLH16+CCysumVGWBM+UiNYtj+
EYBvuXjiv+GRjUQgkLTpzkATYEaGwBv3p6S7ZwKt8H5dpVWva3yUzf7CIQ83TpPB
HaWQe/gsyN8skE17X7dvFGHi5laK/Ehmr5IxYcUEjioAMWZsYFnWAfgB1f6Fddg7
q2XOUkzHNvC9/CJSlBOdqMQmbniDoCIO1zTS2ZlpNrkFDRWUYsbzwK47TqPYu+Et
JST/wo+P5HnUGv/uN2DL3mzjLoh3w90nrJ5yEXgBckD6WwCL7SZcrGFG5CzD+6+p
n36pGC3HmKVTNTRAiTmQRg6L1R1b9+ImCkTk30oXCq6kmXOq2GA2/MAo8301w4/X
Ap01gMc/57vZ58Khnm0PXU3ktTOFDsu7xUl8oayP8KUWsIuytafP9ZMROfVez+00
GFrJmpR3JLG8OxSbLKAzpIxRKYIhRlW6EI9eWHtjmcn58otCYnXq0dkzo4hS4mgG
FZ9gLLdxtov6orUc2d2qZP56CDTS+y3ddmB39b0omJPvoXomEDshIFUi+Lb2Mr3+
xoSR1QMfD8K9Dh+ASaCflCvaJlRZiEYMLbu4oice5/0l74NPZH73ksXcUfZFhgf/
/c0W47N9Vb9sR8Cxzd2fP7vDEcU0UpY45k6OajGsaGxlPM1Mt8K0mJ4xGrZFaC+L
WC5Nvhl31cYIsr/E4YdFOjzCYHqiK7fYI19ATZewxqQQnLh00usRcFC8l0hVSb9n
d94G7qvLRB7HsothL/eEiWUS8QYWLE+eRDko4wcX7vHGdOElksK4lmbmixOAz/gl
I/bIVY+33yg/+cBqSt2njt9McRpXOQddQJPQ6dopp2K12SoxrkYa+wdSa9LmHtHc
gsEoD2ZkYFyAzaXBqBrngzagzhTlKTRiGKn086sNr3PwDhXplqNQcddXbSb+Woh/
hghCY2hyjXUd0A3Cg334qvLYvcfvXISZLMd0Ln3OBFiOeS8ljCq8vBatqvwg3Zvg
DuoZXg+Aucai3sq9kTaaneUkT5Wz9Lb2H5MdxlOznVPSId5iAQ73wP39LWYr5DHx
GVpz49bREuviwDMeCzjPpPsvbWPTha8HYtilC8AxaY0IlZx9vKELRUgw7tPS65u0
hqsNPix7CdHMLqT7IyhssZpxMG0Wp9CFJK2iC3uh+GOG7BbJh4NXLIj2wnatI6Ue
B775UbsWBcYdlOSv1KfiwTGWpnjjUxENuv6D4QJQXbu/usl3aUsIbSsAp3xkPel8
t/MRaElJlos8QLGHtlmnXS7sXDiFgEBzCeDf57qllY4+lW+XF4MLHtAFuHxrZZQt
frIYqKav/e3rTxwoGuAEFyaD7g9eqfngD96IOlc8TEA9j9A+iu/yInDP/rhJ6V+1
ngAkFvgYzprf5lLohrIhHL7sPFSRMeUooUo0Wi2O1N/nJvMU7lRiAVGwIJzr5jhb
09zikBjZKnmWu++4RSSs69owlpAgkGl9G6F9/fYoYMKuyPfyzUMfq9cvsPpZTV3/
IVA0DOM2Bqb/+PfSCYRpY1vnZ1EnAFLFJ2E8vRhdxwlz0IMM+bvjLgCMOynQkOjr
BsNBa25n53ruep1bmHhOUFleF+ctEGkta/xBXa7Lpjp6m9XmeqmRsUlAPFaI1BC2
QK1dd018zzlFQL1ZnBMgnFcAyZ/KWKuRDAdA31aqkqQnK8E4iHeTFRgVqCLMBrQy
z9yvOPcF27CxFu+Ne814/yUxQ+pA8WGaxUvVLBv+TDWOgNc6AXa82Z0qlZ/D4eIu
mdZwJlr/JYhszaJuxCL2e18OWl1AaiPCxcwcaij++VI7maoRTKSBn+FQvuOca+LR
xw1A+IETcR86X4pUZq6lXboWttnmNSjjKVDjEJdno5aVqdUIMcF1RzKKHm4qemU7
4n9C1+vOuCY2rotbV1cF5kY6PifdkFvFkW9klnxBYr+Z10dtgi5tmPrDePI6O6ae
zca+QusMBHzEUzfIz4f2cGy7too2TyVge74IUrwXnqRfWsKwbfTsSf/kzd0LksFX
/UQpalahKkKWAbtYh2TzLzY1C7e9onYgPgPUvlTxy6l+0AqmA4MO+ouClDoZviu1
Oxvdp4/kJb8g1rvi/8Qw9yAtXbNhnxhvf8/7km139hIk/tcn14w4I+Wzc2B1GxaK
v6EFXrzwFP/OUoECw+7gfMjB39KnnLG43tS1uIujax/C3zc8VNg7amuweCmZ5SMT
PTva+UHE6708jJS7mzen4nmAaZJT1FwZQVIjS9HPDd80xT56y1+7T3930dPEgjF1
fb/69YgqoXTFzvyv4caBxXmDGpToiq/WIWuQPYt9LOFbfEHuuKBDIoYvuhDhRPGD
hgTg8HKuz3D7cuhoq48N2o8NsML41WbdapHC8eeFnu7T30OMOq2r2zOfkXB7AG6q
EOYUW2kq3RLtAJuKxxVVVlsf/PMltOycJdD7jIMfePMCgamCe3kDaslHxpBjOYaJ
bi3PTcRdfGuLTLD/xhIj1tgcmi9LpGDDroKZC3XWuqt4cjUtuOFvUkJOGh6dD1ni
BdRz03ypybT9kulPz6UhxA1L8jzVB+4zcbGeXWbdXiD1NKSYbwxdccvC3GvFe/+e
uVDe4l5Qug6pk7I7GKUi5vNeNT+BAHivrXKjNWp3IqLcPOhb11FfogwHwa0HCCIO
AJwlVsPdrJwSmaNRbG3wx5XQ/6EHCNR8D3CtFGtzqcWT8fLyZa6lxPxeGWXLXSrQ
2BeEL5kBtJRnZf6Q8P3oXlhC1ZkB1ANPcBEyLszP0y7/HxPW30SYETjwqhz1WydU
sYGojuCeCz2S18WgrqVyglQx+keE/7+CJpOGNNRSf0dM9U6OYjgQHdtTj+pzVxuI
YweW/GKK+R7wUnH5Cc2J9kS8o1WcDnZIYr2jX/dXCZw4qMNdBD768nanueXELZ4t
85SJtR7ZmsMs4KRBDAT+HckO8wPxjxBIgSxcTKj/hvasiCyeM2ml3hnbkc35QmBn
hji6JWiQN81CQ9Yu5/iSazVxs4DmeK1Lxm6BWLW2u8h3iejk0bi5Fd+LzRcw/2Ot
TZ8FwkOrOVIHH7ZHxH+2jSbrIF/K6SI4J0j61x0++w84zEe2/GjWXAEhvMVIpnxa
jriSnhqyFzWvSVDChZvIGw+gsfLEw7U6rWkb+CFtJBWVDJ+UJiqKVt2SqxkMBcN6
6Em1fcElIc3j0vblXWO70NQO94dgucLTAxjWfauIqYVbvlHifJvPvLyBbeVGp35a
jhHuKyCNmY1kMQO16vAnZWDcuxMreI0ggROU2DT6YW+42t9v43XxsV3NQkcODI4D
sFHUpCtegHxqqsDazlfuyk9r0PNNMguU3hlsh/px/UefH1Ug4IVnOIhSzmHgyM6E
XJ5afuRUglTj71pUPz9r5T4hVfTosbH15lovD6pbpsUfVL5jT2XZWvo+exUfMttb
lEX73ffWdYiANmYGDVRDt+lb8ihAoyeKc/kLDEC5gpwobwrZRa3V9cHVVqq4QtQj
rE0WquGo3v4GIUv/dXlZT7hLJMMctWFrC5j6C9VPkUKBfAf8Xu6ljk1dsQWs6xI8
B7EdFfv2H28SSF2b0uDODOImfDswguDTJoF1/iAjsEOicl+e9P4TkxBzzz7dFGCq
t7LFGbPvhsBmJFIrQiW27EXaeH6GTJ2C0e4EaCCVnWWFuhv7mZKHGEuu2oW8Fo5N
8SdnnazVIL8y0hmsgSq4oqo434Kq3kaTddVrUvTSvmEuakG90Am4llqpmJpsv6rj
29361GfrxRJNcQegAafvrHMXq08HNIOlphbQ+K/rtCHY8SN4N/BAbMPTHGu7PhQx
+1ukKsM3quGrPQ/o/EfGWahKX3myZCtefpjHAo9+Av0bc4h7/CBfo/s6LwPwtoov
XSkLA84W22ZoFJdLGXfyUvUXIba51ItKROeTiUPSw2TZ/+OxVwNNlXvgn16lpQ4l
02nYOYdDI//KCS9YW9zEdMqsfQPD5kYsuoqIfDBtVhuWNwM41LbPwFNBmowq56ww
JMJrwcUYsKaXWl3ix0m2PfuW05c4jEZ8h3htcvQY6sgpuf86pMDgN8LSbSi7Z4pJ
YuhTGQXLiS2Jn3cDg5V/KjSZ8ZTsO2hOO+HFaICdUzFpslNaKe+11wQjjRa0Eu5i
lopsMHGw39jQo+Tv29ze+5LqF0mkW0hr6+sIfM5PY5rojNCv/8v+44rA/lBx539v
aLhWB5IGDOZTCnbTXyVnJDBcHFRxZOXXlPMusHCVjl4VdmRRhJ+6+v7tcKMI/wqL
D3z2jIgGdc2ooQEB7NAZgAlqIv2O+aEGE/nS4ifbhQggcvX18cgJSll+LYdDscVU
vrpIq7oGWnbmxiTH+HLodFfvFU4c3d5MSlTg994elRzc4RNck8ENHQLeNLRy8ugi
5f+tgGaz9X9c/rv2tJHev99PLoTMQmgLXLdJ0YSpli3mHDEgbfEVFlR0pChVLOie
pNX4ZnXvXFIXD3cSWV9CdvrV1yc1OevflBDOR8Ta7NERPk1Zwrt4DKsjdjvi26La
6xxTOoipDU3b3tyWuFDo8WXM+I3qtHrDuPo4n7+DdRHDhYdd4RGfY0BXRJkcMCp6
oCeEtZB8HC988X2oh9bddM00H6Le+MuThxKBSIBFqpODFNr0cN8kFCeLT/CkhnR9
bpSqu5T6OdyF47jgn1hB0qpn8ljyIWyXLuYLGpnH4/5mScEKhVrYr16PMpj8Qs0B
KsdG30ekJCwRcC8CXfTfbcGjltAmH5HFk0+D6gyg3UkVZVlwR3z6oQSYL4i8nEcs
prEH4V/xVHo37hhWlHDVaAdhwp75328jb1EJvh4QXhjrTtIgIenmCEVQjNsMrXaD
5xBB5g46e14Tv+nUwiUIpeavKpXYXCgafPtt74FdsXVU2RsAq6e9m6DtBZVKU0/y
p3ZDNOnuzFOqYq5H2Bt3YCl/3CpjlMURg3ndVt7EWMOvUafUh3devU46IlYUBs80
PjZYu28hD9q6Fbk+B7/NAn7JlABfWd6Oj6o/Z+9T1DlODARm767/MJuU0rkqh85B
qy3tIYBDI3eWDPALdfIlUH+yhxfDmB1Qf5csnysZQbAXv3zl6valIBB/UDYTXKp1
DrwmyR2Il2GG+vJosPYzfKE0IVfWFzIkvjkEIxjD0zFbJIgACmDynEChO28Z6Hy1
WnyRi4aUykUjbvvY2F0Bsbwsp2fn3/RD9XRJYDIptycvbOmnNrl69tPSXmbTO96I
A9Z/HPkID+ityCBwU4iM4vjVbpWOPmC4qxdR2T+/N3gZqvUnIbB+yJU00AzAf4Au
PDRRwf9+BNP8BC0TteW2JAdl1i+WlQsLU1LVMMkFsQmkDi5OvxVA40DDHulK7XTW
0TpwNopUoGsa8Vsj5lCKAW6IQTWhyoOLXUeXfA9eDGyhSXflfGVAvwVqAw4Xjism
8C0D6T3vT2b1mocd1tcNPZZIIfIYoTgB4tnn00cfrjrGX7pc82eZihXiojwdajcq
iST9EqdnxNs+DL/vQjg2cqp9xQur5V3uGqW6F1v2Ebcji885XWV+0L+KTAHxBdeQ
Aci+mZDGI9xxEWKQeNcWBxW/KMkvDXH2M47yRTFM0vr4b/NAMunc0ZNZmb2TvkFs
L2dwWz/FEhyPIGXtCZd38Mhfz+diQERYU7tCXLM+lzWRWTDP20LvgJq4IujzpFZ6
9UnQHlLOlDEstcFaTptwNXkJkOfsGpL8bqOhE1eSPEr1r+GjxZg68TBkfWNJNt6W
UX7Ya+oufCjawBpE2rqe/6AwvyMHNtLQgUyHFDHCC6o4vSKDubIlGgW0SLcEbBTh
86vkzf4cQT/USotH8sQIi5HHRt3S0bijgoIzluRG+bpNGjXdXHpsz/An7Yc0ilrI
CPFq5RIp4BSAin5I4gCtXrQttENxw7Y++WcyTrtciTxdbtCPgedJXlAbu9L1/Fwx
eWpB/CfaGMbYnA2zZURc9XjcGh+8El2bSyTyhLB6OefkzhBN/BAOlUQ3Mb7KfaEs
hNTlMGOsu9OPYKX2b7ANoLFsIiPcBwxCAnX+UO7ztpj2uyjwsBd9qacCptDkbiUd
NHEwGl4P3Mr+4FIaz4oGIqkn700C9+dTBkeV+l321m+3C/Vee2pXVeA2a+1jIpvu
ciHtxgwKHTyhqCPOwqZm4JIRlkObL45T398S6xFnsin7w0dCfmwHEp8SSvDT3K+8
XmNtQg3zYgWkFwTawTEkDwqm6Mjq2ffr71KqBD5VS2fJ3UWlMfejfV2udW6bAxnt
hTVsYMX9MB5oBei8Q4OUNn+N2AIAm7bZNQr9lIcLRsVhUAUVHPlInDDfK+BF/05r
uaoRCEOGSaeRGjmKn03BjS5sANL09ssDcgw2XpWE9SKiM2ozS+MjPVrFq4FI9NIy
vcAUi+J6/TqidP4NQHQvmRho/1FyiuKIzJXdPeTP/zTKGZROj7DTlcSgiy7FpuqU
uPvYZIB7Xb1mmDcxJsou34TG0PotYOs9lwLxMwUXewtjJVf4e1Q9scuQ0IoNjwlM
EVilJR9Sai9bRIM5nJ4S6HNl4zVKlhvMNqnV6GNYufyKjA0dTFCpYcVB1AvWPZMu
SXHkeGOaIlfalEEp6UBJy+JNfcOY74qWYo0YPYuOaR8TAD9PXWriSaB8blYoIU4K
hVyqgSmFSlIKqpSc8/V8TmfC+iSx3Y5nOHDxOJtBl2fbI8CdZ5XlvngKjmgIk5dS
fQyHVW/sU0IBJQ5DO2hIJwt1yF/ol+a9bmuURIKfaOIPoC4dcI9A0wSE9GDKVQ4A
D0fhj8hKhkwjjmKdBOG1WPgSHapIlWhEdaOB5vZcILVUkjThFiCUTGr/zNd7rgs2
nFdgp2X365CfEiIiMRMrsF0GZ99F6/RaLV5e7A2TShf8BvYwJRruYfP4uh4qJa6V
PMmDAT2K3wTT0TDwIdTr6ey8OWDwJtBny1K4fwjDjsWdS1iEN+K9DpaKceQB0Zqk
IpEqvXgPF0YGMIFZJUmguVPnhKVgAt/AMkEhHAapeGu7QFxUgQQxt6J6f+9tDakI
2iYkBuvE+fTMYNzaIHVbHP7O5QC8kuwcI2cHBUD5hez1uk6kqIP4Kzp0Q7e7CZPn
QjmgJIuXJzMMagp0g8jP79TfyTLfkH88NluwzIxqicZXhyFQU9HXZDf+KMKhMSaA
XxZvAIzE3boUNYrPn+P5yLOcWtQ3wgarQAQhgP8QiHGflROXhMygXNaJEO6S9t9d
IKETxVV/y0K7j/X9TbX3sq9lYSF7Z3Xjnt5VyB/ULZ+WcNrwiBc8/Z3wMps2ejSu
MVd/mNCjC7s3fB3PsxhfYpNYrCODs5aehTH6+BC6XDqKN+qHsCf2xBVOY45EdwEW
1sFepFwXl+lsjgDWsYYsmvM9NByrxgo+QQ0twxagEa9RtBdDrVLrEvijFNtfwHQp
LV0l+10q0T+xhqdkXzztrDBsy0k7Ri5K396QC+7qTZ3WPqe7ZBoxhKRhk3t3yA6M
hqDbEIvZJNhoWtCIe25C2dVQZOwm+p2+mA9ULZomWNLN3WhoJDdPXBG0aTA/BYv9
VAHYy7r+xvGd9QIhv+dN8Ljj9sFvc7uiWx1O6DImqHj9TrDcoAyA/KgDJo+0189A
SdvFf5CLG9bCpBjLZ85dNKgl2a1Gmu3TaKur/0kiLhnlBXSbWiQx5OoxN4aEaaoI
Bq5af2YYO8kIAObew+tAnbDyDLLQWQrnhEVlD6/0kP3zcP8UJ/20rrUR5e2jr2pq
QMGIzgE9vBUj1qiB7nx7bihwrnmVwHQQuo0XqWrvgsLUy9nJeqy0djxGH2nMONWQ
urkHKLuiy4M/zNzNzLv4CQM/QGLQ/efZh1O4YAb6aPReuOhWpkTSXnDQHcgQdH6a
LhChLXODZxzl6Az92VTHEFvICZWdIz0hLaWoJ4NV0QGukcidNi1WbchyhMpCOZOM
CA62uGEal7qrMGi9C4pSYt8i0rcJBN5owEA/pPyKMZlxeZX8dmySTYp4RzrEKDU5
0XaV+6Zv+2gjlfMbh4qjJQyLKPUsI1VtLxOt04327EymBTDtPs8gqGdqC/8hcGlA
OfEwseUjClBEyBZYZ0aEbydedvJPNlBV+XunaYND3iqCFRIuQ89qEnPYkTTbpMQv
rwGNhG04WZyDo/Nru2JvWGn+gzUa9TcyUqsvorfylLAH5CDHDPzp9vWehSEZrJgP
KlACifMuisSV0LAV06cI9Hz8vfnxka1qJ/lFIiY4HF0vuI7j4OLLJXUWDs2vcxnh
duuZNaRz9FimNAEukPuN6BQ4UATGu1Qnw9ztThDChBpQo+qjwhEDYfkO9c6GrO4F
2nm7DiPNGowvv0E3I2l8yXTAHf+5vhgTeXrkCpEQ413n9x6AXGJwXqcukG5OoXXX
Ezd8U29JiwiNqqvU1V0CEguuGbT/xBXJPVOJYMeSLXt6wob5gjdrPzwq0uknhhYn
h4DU8CTUakFEBE9Qj+vnTY2GhQkL4AvHZqDY9mxVclFQ+RtDuwuDB8bo3Tx93A1Y
mvm28RZFQ3nNma/WJ3bPjBoJMvcnQlnNrF6NIl3A0jgIvQH/3H2UETKW2es4oLDF
UCtXiC5av43doCw/uc0q4aWAAWY2cfxa3ixiHpwDfgSVnv5H65BrsHK6ppYQxwXg
+22AtnXXcSV0ZDzegJFyl1X9xSnye1sx5pqKOEhxkAylEbjJCh06lVK56ehgdCnv
7v6nz05FeJtpIuXtGsxMrld+kgBAZskDgmR1undG6piiBLkpKb9DkNyHWlbPBBzs
E9aCZsx2yFxPkMuVm3OtlwCWkT8VfwKRkXjvOzDx4Q3V5GwxF+YEmNy8IE7VmIEY
9GrxAHUe3LxnGKtzD7D650jCCluaw9tgAiqBl2TjGhRjih+LrHE99CgCk5k5HN4n
dRepRnev6f3H+yt2IJ/VOHPjQABFw+ii1woigrpx4TqCEpGI9Hg/9TJOWeww+j7L
laQbatzlQcVttM6zKgY5kPCzFPJJM199xNxxRsCZBAYEKF32wnrvJpt3PwNloEgb
Z1NM0NDNT3AZClCVXCjGIZyVDi947MjhhNAlx8evpDuWXPV1xfO9iWqmMpx3Mn/I
5c5a8blffUBEGKsqZJ+G24nqfE5FQw8+YYbKPpey3HOIe9GVOpGm+agfxZ32BNaw
GOlH1RFLH3gLPmjvqlROnapAHQmivXfDgZvM2u3Ux2iuNbJDNdbE4ALL6TTZibFP
Ccx697wDCoXzsMkYQSnT5boAWUWr4KuytWJrh73F9G5wBFDdAlAc0CF8lBD3W0ii
QI3UXyrEqjehQIvwcCV59GxUVXcwyzgcmXe+ogH/J6s2sRV3EwvH9Xi/wjyzqLLU
8Xdm24sMIKwhIXQzi6OtmGuP2HXKLTZKgYftpEQSJzhm6MIurg+y/uL3B/HRnNPx
7z/6kWOp2QP+RrfiuTuy/NGN9jBQcotoRcuKkX8UgESP/3r/JOdxx7z1kH9Dsyf/
JYsB9+8TBIogdiWpwLoI1yQ94X1Gy51FI+ucL2IUlWnzy4x2oj0BrROcy8Wqah2R
Oze1l/Jx6EH4+fQyohwrfQwCQcx2Ru1wr1PPDlHu66EQ3KJh2JQ+D4HmHQ2lnmdM
w4bEIrlnxQ6zOS1uaXSWSxOioR4jLqMdAxWy0TRCjfv8VFbm20Ao/ZBzvllAuggc
bG20ItbUThgNcUfrscQa/jvk7bjdGnPJVVMr+Xr/8srv/ngNKiY5ZN7GtasS3lN5
PXAQjkogDVY54si4ULPfVf3jvNUSGA4+lHD9XIRbMC0DXbubQ1025xLIOIYetxz9
05ffLALW+vhHO/ntriYYB3xwJKGfSBkEgs9fMngAv78p9HhF5Ol7/7jY5F8GXNbi
BiBxj4CJDzpz59YbtE5ia4DhESWSE0G9iloV9iMzB8SaTi3IDJe+Zh6kQmgI4543
MTRS9aYJ1XEpTcB3TFsRO881p3R4rM9Ew/qiiMgl1A3QzIMjguo65v+g/jD5ZyPF
tVQLEHxuA37npSeCKB4d0GYvWuSpAtj0Oh3G4bYIDlPzLSWklWmt0sXK/S6r4uY2
4HFv6+Hc40qIiNkeRuGQG+eijvGGd3l+iBlkKWlVf6Up+mgYawwZPN+OpXnKEDw6
Z/8ctB7xaqueKJ87IHaeOD7yDTd0HxoBZJuS1AV4kHoPRTDFJck8vvKvc1/AJTiq
d7EWL7uLctq+pLzf7+gdf42taEt0XaHCyDgc0lxYQ/9ZX6QcXyehZGLnss8yycsF
saBgDxHQXXbRXQwLWkrNH2cF40OeelnsTzpX4B8oLPTP/HfpOF+dx2PZNaYxKXVP
jncWB4X6lhlc76klcoJhUxxz82moe6vjbgGg+IA+DR4tflrvBnoRMO4r5QkxwJxR
jFRZHIHSnvGgHbHtDHpApcjPMOebS0aOqDe5+WWJpZEp6L8SVOCw4m5WNBNSffkq
mJBsI4k4lTVXhBgNSsv1rgSlS8UVq+yMjnGROZaEDqjIWhelIv0dAao+eTBxwXg9
7P9v7tnOk5sEj7F0wVMvXpjT65EyO2dHHuZUVykJHxWow3+RFPf0WzHJbnZJG8YU
UEQjqFJBxJ7AdWkGsYJXL03JLmOvhu6y6qBpF/BQFQPxTiZeKBt5WnEIPBpZkJPF
DGsBtwe9nwM4DspzFY+sQI8InB7qlPq2tz0zOWEqI3s8jBp/29X1SbaRT1wNSy6A
qBaTganJxFZNd0d6YYiS7+EPm+M1S377oUlDC0AjXb+wYZ8IYYXjz0yj5Plo3m3X
LB9Tvr2i5T/kly4WvjyV/ZNDy4ZLFoIsBB+99lHaZ17v6oSAtaeeWL4adt98x1aV
ssMX1axsNdS8omXEYrcUGpv+/FQGoWw+oWUxuH8aqhGeglNlwmYTe9IKsPyzZ0jL
OGYNv8M01UbQ5QsjcikA1Z9JRnudrrjWApj4x0cLxKQykNI7gnO9vGCOEhw3fuGM
wj342V0F/hNvyY08hb4IYCr2ewXlF7JtD5QU18NUzM09AS1A0VHNYOrvnyIZsPdu
y5zti4yort6FZ+TswU4E7rty9IH/1SpG2CZm6FkJSx3EKaMb5TZkMy6rQDsRskmd
9vtIRX51aNUESLJpbstQzez3po7o1/0AziDpCLmBGwYxuTomJrgFgBLGF5p0IhBZ
P84/qJyG4V5QdqO7KsPqcTCdhB+izVGwkNjA95JAtxcdGp1TeGRicOBwCWxR+Fq4
0REDKNtUCL/+5H5ZOhk6utTEd7Yk0fwwb8skGA+YXXBZ7T2o9+fqQkFgLspF4ZZQ
pwuK0F48dn1VBqlNEVQmaZxUFB7FJKsyO9zzQCjrTXPfEXpUmfq09bF3o37bu62S
NFwuj9FHRHxKGxoUM30IOzwCagmYm0MwLyzKAUX2pAclJVccLvBu/cqxXwh0ro/W
yvxghd2XXa+E/CmB7LUM+Mq5BZRmS1z982T7ZJUpMPygYY08jAYuNcx9pmoLqCvm
+CbBnPeX7jq7OGV5ySaZ621oGLQpRTYLMc+O31+AT4L+S+DMdpZJtdPjAaljDaM3
UnmGuy0+CFj2GNJk0lBu9Wf5bLboa/jiWbdBknVEIbXy5zqiuh+sb58mPk+eu3p4
Mm03G5D3wLhpZerOrADKp9IetYGBzsE1Q+wxJalKXGbBegn9DPNNxv9JZ9Mtlb3j
9Bhz6ZdPATt+fEB+ccWS541iwsvvxjYqY2tL6vfaYh66y44YcBBF6FFV8AmDrFMp
U5SM9xK+oOowImUIyqN8O9gm4NEf+jS5bJ9LYzo98cnXChyF0whxzdMGtEmsymNI
euSZPZnJIBFlJSzmaVj8pPGLRm6oZq6rpYw/K14JPhvQfdGxuxdALQ8bT9z3BwUv
ROxaO6GoVYhy67tlkDHC616RTGXDuE9rIX/LX+kFExPZUhFuPKmmDUfMVXCXq9h5
BEW6LYJg2gnTrbEewMIiY5tcGggxTsALnGcCy6rV7tL/bSne1hTIbHjWli40yn5W
dWDFHhQ4p19JDuxV6BQS3+6XkU+11Ym4OX2m2VBocicorQ95XF8B1XIlhTl6dXdm
jZXpoTs7osu+4PyaH06WCZnEF6FzBnDj3W2fIb4SCFj0OQIeuYMVt2ULQcRqF9G3
n69tHxVR9BdwKKx8bkMkrFOJgqPyNGDSm3Qx/4W+vjL3x9Q8Kpv76oV8z5EUQDEU
u0JEayK5mfe8B14yuYos4558Bxl+rWdlbjqx460k8GULAeVkYARoQOkGiI6OuwM+
yE4x+WEzy8Dmc47SZcJa/SYNDVxPBo3eMiTzIvC6gBAoBGH2BEh/Zel0G9cnhbKc
Dxwpdldi4QYQbKs9MUWyVdhMDWw6aQe6+OktfbyIItvW0lvhXw8ecsLuLrfqg0CC
jpRAXWj6Fw2G8P3s/6/zZjmracXGKjeYrGzcos5yKnH6EwFBItr0t3+lC1MQ3Df2
HT67DWho+T379vcSostJQ4a3g0TKOUXoC8shyQMjvS99kk2DFCsfkExJzV8H36rp
Cg4x7/MJI+6af+tbbJYIV1xnV6Yfjbq94i9QZVjgZ5FZK0J+t1TO/GjY/JiQqitw
H1zJwYlvo/pIuFM7VL9jIB8zE9ajFi51aa3OjMtXf7+9BdmOF0HZ8H2gSCHes984
sKvI29yOMWtEvRU7DiS7c/I8Se3bcvVPLulgbacTNAbhia4FwLpcRQoJVlEMFHAm
3unkNTruwdyUomMriXy6aclRz/IW0fx6Z9UwmbjB2T3RQ5nCgANSxHMddM1P3Zg0
UEtPmMNZC1Ome1Anoc/czRSERIU1UV6MFa/Dth8YQaR4TiGosQdYkJDi33iDxOxb
AD6oCEXZGos9TBlEPmTa6I2hhQ4iFI03zjFwofnfko/QXoZytctZ78H9r8OC7iRr
TNNbaZ4CFcnm9Hn5NjC7xWqt0E3xytia4whLOfb6hg4MOsg6Ra3OW4VoGHLhoHIn
iN2d1ewCFc/z29Somvq7OBGyxtBFgszfAydYgtxfFrKO/vkRaOh9CB6sNnsQPfUi
Yb2jVf9CUOloFZFd6ChDCYGSGXCcmq2+nxgKzPVzj25ur1DfLFV0I4kiWmkPJNBZ
Atb6uljYTzGgeg7uBdMBXlumjX2KtveIT0ph9iqEzMsvuFJn5R5zbgPnnyqbvX8g
WL0QUFB1ugOlsqnJgco0tYofILQTlSff32UJWSc8AwGUib6Dcp1LP2NLQpyHeWex
mL7PTknRdiiG8SCahd19P97SryiRbqexg7xS8tCy/tb5f77wY3SgANwKfM8QvunH
VMA9sdM2oacgD3G5t70fxohehiEIWg37H3vZjh2utmRYTZmSlanrXRi2kxTnDXlL
S/LCc57IBmsgndsnTJ4d4Jqaj4J2Jqb1wYJ0CKo2PD6lG2q6Mb4zAoISbEgg7pdX
koiXyA1p43IyOzPhzF3Fx8oci3MQuc/7Xr9P6M37acibs9TiHMj/5qY5CnbdTktS
BZsAzhduu8v2Fn/qwjfm1+ysUD/3wuMlWbEb2Aj2k8eO1P53ORtZ1vC3836ywwcs
m3/58X9W1+51SIke7CK0mwFBFi7VTmd2OqMfVJRX8trBgoDjyXL20iIADjmNfu0X
ZvNCGQTKWWopEErNnJ7JjpMyU6sBPIpKKnjxh9ZUA6hclUdSjag30LINf4OvH2lt
4kcCAM5w5xpofiDVBRFDl/XCOnPEGBFKsYRTgj0kZvKYnfZkYsbS1O49Ao8Y9Mcr
J12eVzAMTFJluAp33oRZSrqo7S79Tie9kjHuVhcmarjFwIDaZP6nXLOjnGvR4ft1
HYVgmiAWbuXfIPaDG5oZVUGvDv1JR6Ag2861KKs7JGlk0FtK2aTxEJF7LtJLQOwK
OZXM+mfjnPNAedOT1ltu50KGYkPROIyRMHzvrk0sJbEOWUPIEjulvB9fbUbk+u5e
0zqVnfHviUfTKND3LfPK/IglbgXiQ6gE3RfRBnnDc8WGeFUkq2Gd4gDM3B5s5WAR
pI5yRg8nAG+sf1MSdUBwaizhA4ao15btmtzws/G5pRmh+bEA2PIYxLtj8Snw1GiW
M2CdsPYunIn0QUEySqSH2MDXI0NGFSt4JJbsqPa42f3c0JkVLbgO8IxuB9l962JW
Wr2v0mQE0Pm2UCdfvTKBhcmcrbgQjFeHht/t6nllOfWiaqchagUtQvDngu6kiR0U
eNQlhywYj/LhxpSi7TPQA5eYFYgzZly3pJippCAr0016J3NUeoFyTzTzVzpLVUfA
BtqYTE8/ZxLl14N9dl/XoZY+C0/nrOvzenK0Ku2C+NluEjL0UcnbuybnUt1jeTpO
o14U5Mz/GCPWODq9JMKtpFVCC/0GyKoTBKCNZN36GYg2CxmdixbqfFubHQIwZaG9
nmSQIRuw0D6SpmKU5tKoH87go8Zy0w+Nyc3HLUnuaJgKC9EX5T/NNoGeUBduP8Lb
yezOaSdYmoDxi1PRD+UosN3m86D1i/ReDDK4SoQNXlVWO3nhuayyQTRSmCN+MOdg
tdnPAQUbiZrPZ6nK9qk22f3Y+oX1ofG4vyXl04oe0iIAlK3VuBPc1Omvp75ppSaR
pLekT7gw50FSoMFxTvj+Wz9WdNjGuBzRd/rWV51KYUlYuuc0FELMsdm8ta1zPg3N
ik//3vH7SjOjDtZEtZeVm5TS8q7rOWxVO2cF8yFOA4tzxF0ZX3INiKyEEpjlosv1
93gFmPzNrWXgCvqWckXLB/MEx59JDvastTzKfiBYHI87LDk5QXBxGJFfeFgWfJYP
LgubuNQveGsOfFHyad8PxtGqDr8/D6OtgnwhLroEo17KUN8+mE3fMgamxeZtE5qn
9Q9ypTXPCTGaXT6zRup2uXLTqjtz3zNieUrnxruJqsAdzhg9j0vVGkNYHE0sr5Ji
EfYcbpnX8J/HDN2Ws5tctDV6rFY26cgiU5YkXPYe/mexNMGORQlJajmNuItr+2Ow
BLItgyDxJWAsv8zDAkbGQNzZ5omqlFfjawy+5bG0cq3la1ZYmGetIQMosBN96Frr
+8OSjQuqHsqejU424byrFgImhE8BXuGeCSjlI40HCbjntsHhAHJwhcrOW/8CoLMn
h/O89ZqthRf6WVUgqTA+r4MnqpPOwK4Bn7WhUQavVvKT8+yUa+BuMj9ANs5cYdZt
dAd0Q4gNHFBzNbwaTL/jwCZrg4Ay1IjGWRb88KxfcjgKrQiDgTqJRp445GiTvw3g
oAeF6yNchvivUTkimrOltXgEsg+lgxjhIzsfzWDCSQbtRjcCjtDV6zJuOi0lT7EN
WWgq7I5H3xSyJ7Fklej8bDaodflLKyKwRbSjbziw3rtsARTL5iItLdiiFCzVks6f
tEW5/is6w0GfSUPHf8HDD8EijnfaPaeQ4cUNsMsM+KSS84NIoI/q9UVYIYQgdAof
HJw3zn5rXctfRY0R2z/VAkyGDuKZFbI0NJSwBKxMs1k6EOxpyvaFgQDpGY2+ObsV
U3/2T07OlRbs//o4xfmS4B5B1k1a5yJaLJbn43m0TsCXt7Z4IahGLDyAUqtaEqWO
R9HHtoEl2J/wamkImA75P7OCF5CQ3gY52UUD3T+3zk7zhz3OFewFZGqCl/wql0da
kf/Pp+2oHGLfIoVL7JbkoeVQFghLdeM8OejWHVNz3pESCardPF7/byhIDN1xk1km
BKNs5yFWjunRYBh5qRgJz4Cdeeg6aGL87ItF59AUX0AS3l9Abm1s6cJX/aoNcHa6
zZOT5UcUiVstrtpnIu0WYo0xtND+G0WmC9f9UGmUWVgTMGKZRiHVhHeQpTGXFT0G
aDid8RfJQghNV1sqpYLbyjnu7QMmcprwPJlhOUjG7l/zb3bkPWVM4jsHUjkXd75u
ozi7h1z+M5GSXa1OKc4tqav5X5va0IIcuDR0/Nc6VaKXEyLB1ffak8mJGRiw4rEX
2DbrL7UYRnbEHAHtvCak4aOAqSGxZeZwyhMYjClzgCuYVV+9MFkzkns2wsZmr4p0
PSkzmhtGdj0lYbtdOcFutfmUH/7pRhe6+GY5uzrV6ocS9OfLtNemiW2kHKjWHopn
h2tzAGOiDABs5AfNiK7r9PctNh4aiLA89r5iNac+ECmQ4NjXqgnM2+L6yAcvzyji
nI6VQpNFHOaAz114rK+J7bX5LrBlx1tclnVrmxUlU8F7hr1ZTdW6GiZtitrxMzUW
/dEo3ZqHjUiNnjw74XZuD5/GWkAfNcWudw3j/zYKvrPnhtGs7vIfKqGjVohXmNdj
a/IvACVrCDfQrdPlJnP3DgXsySId2+IPgo/6/xNSvz1Y63j/LEEcHq6eDIAnp9ja
PB9YkzX1z79LNTfeoXwS18agr5JfpEjr4Sp0h5Mt1ja996hr7TcT0OcjYvOFQ4Db
dfHOk9WNgPkr4pk584YS7fRrbXzHhoJR5MrZ5rRpnlos9ye7bKLGPs1UCDsuIUAo
Y1WDTZiF9OdwCAvGqkf0aIAJGJXEawIxkoj3o4V6i1KrIxG9tbMMA4GwenDFI1Ce
QZPKMeQG1B8JFxTRB8lWKa7FDnADnsywhcVPngDyWoxbBwmWpaQmwPQB/HgtOkFj
n+JYCCnlUA81jqa5zeI/yeO5EUurgKN+Be6lTE2NqP4ma50HlTi4GPQHgoKEcMoE
AtFLp7sgeKX+FpujlwA0l686Emth+mKGYVC0f0e3TA2U+wYMfYXyd6mXdWQWvC/q
g7gJOBWO53xtWJ+Zfoj93FYVDZThH/eBN179n3Q2ORapV+4Or/sW2EJPqwxCtE+6
O0zQytHE4isJiJXG2crCDqmqrrphjrVhJgEXxZYPbbf3ZlrOjJim1bU7Ona6KyVV
7TTsmAhPHR8A/ppd0HH5M89nk00mwoJfJPRH68AhHHCC6rAF+3O9+43M6IMB3+8A
yU4HnK6YsYDcM1LZ7tPREWS50LXhx8dAvAmLnlLRp9xGmML5apFNUA8HLwvHYuck
L6xLDp0j1DiH50sAb4+E+0jGgpTSRy4ro1tKVpSF4wuTeCt+q1t/xGc1DFWFl+DO
Km5lkoiqka66Vu5RRQ6fJs6CnZh5dNEdTIgCqcdZcAXwNqyX5qumd4fjS5owfIAg
s70AtIVStId1JCv5gDoojkgu65KuH6I0TrUnQWS0+JcUW9i5dbFeChHesI+QsWMg
G93sddFvPGJ/nrR9SKLz0bOyEsarP3F2ItY9gcTTnC5itle8dYweSH4rg8fNnX6m
JvIeCstemeNE6folSnhHjHKSrwS23Gus72G0uw/+/wVnCPa2zENUM+OEgb7FWa93
pUj0mbvRpgAbH2WQvCw6Nh3oVbCOAWjrRJu1rXvfD4ZGbg9GISeiW2W0i1Cfhya0
hFKypvF/U3Q151All1kqQfatFEAi8Xu9lL9PIBN89Kc0ByOHw6Y4UZyS0RTqp8TR
RGnaQqnmZfUSwJSKwB+2MOVkdsnk2xQgwS93AQG14CSGn+3Ev86b5uhRvDumjw+l
iPtSXk2Hd3NZAHaGT/py9zj8Ty1g4UB3RupdDM9LbyjuH0aqlejpWSn6lDoOHX1f
1QP2jAnnjE6UALuRqszDfMBFeu8fp9KE3VV7mI+SDI58hUkPzyesNU+ChenzKT/e
ng5orsdQG1Ya9KI7Qsr0Z40JlPfH8mO1/+xuF43O3SWBmo4lcWi6d9+xS/a2Q04j
QnXYF1m8/f+cwC8YPyKlJd5F2RL7spj2rz+Lv6/Jo8G/empOV3aUNFfIHKYoTHm5
8fKN96hBpPqVIbFIHk7ZpZ3/5KOTGiT2sPFdtGiBwnGpG0xhJOsu2pQKx+If4e5n
3k71BG6jXNjxe/n0KMIywdd2AjHaH4lH6sNBWkrrlB5OQpc0MQNmsfiv8ARuMLMq
kIYzqEJCVOe/g14wQ8ZWPR38vPFwd3te7hagfPhzRd0COMVgaPimEvrULy1zB9Mo
RKM85KPbiBjblZu6P1KHFI+PHmKLe+zzDm/O9pUJUHxS065q6f1PnozSZFMcg5p7
dgrDsW1JKxNVQCD9ePxlLtRzolclTIDRYabzjZPq5Z+5Iu39/IkM9GAjz64oXYjr
S1JLTaTrt4G1beSdqiYCY28/QtY5hIkYY+FmEIjqZx3OzfGEEIUGZPOwZ3SD/Dkv
4P7kAQeOscLdKaKJk/gVb6aH9bwmbqEFZ+H/9cBF1hB5gqAycEpScDZVBqk7F8wL
wLVEVo2zx1ezy4s/vzAZ0HLdNJLaH+EWpH/rMlAbEsyg3frYR+Pj16j0iNsONrdL
sp6aV3AFj/qk2rwAGJk+Yj9XNmnX5kUQVFjUUmsR2NvDBUDPFSfWXBtzVuM3tne/
/R3ZaoaYwJYUN01OyWwgC93ioqcD6/hspZyFnAgGMrFBgg6OCcptblW/JoWMF/nu
tIFEhs0MzAdrt/STbTX1e311YSw7Ol2QFRUEXz3gL8yHNUXkUqapqQYzYrkyTfsq
f0ZyoFEjn3NScCMufRnZsqflJ2XeE/MPjLVsDdlzvJx1Q/v7EtwX6SqQXLQVdRUn
IjF6l+u3kWZ7u6j5jVQ5WxBc6I7a/ly2ra/MidNCdikimkyVL+laALX+DtIhpniy
r1wxNI2kHjJLgO32ygZlcB+mpYJFJjKxfeyfanTHkzJqttUeHGGHvpvwLedNIx61
L06YcVBBGUt0s77azLkVRVKzewXQUNu7vZ69ZgrPODy7qLntZ1mf0yCoD6jnfvia
okGg/2MIBwr0r9TNeD1lr6YljnGXLdId3ONOATKN3k0uOKA3QbpMx7PsKbB7kXJr
rUrdJBFHryDiXlbvEfxxQU7wutxBqIxyIS446cRO99UD8bwWEdEqkT2Hm0/9gnjx
OxuY9H7mbTRj8kHw2Jb+DABZISM+z1ig9Y7zLLI67922ddYmLahkLcwqUcfG+T/2
ryKicrqU47uuwzc8rAmy3cCWa+Wx5+x++46KP8ykoxaYbXYKoTE5MI5BryKIaHcr
YPiiCe1NAYKBHwfrU+Yrp0GBynVvvDCyqCnpvpuFzrx2bbwD/RmuKqkPCTvY+R1V
3KhYdcihSXnuJic5F5SoEEjZBtg6BYA3qRdNdaZw7aCdPn9TezQtzCvg1nEiJHJV
gZXtXP+qDTiYlGH+cuqcM8dp8CGD1IvQQ/J+hWwgO+lsGfvlQ+P9GGCaUSjl4/Sb
dPOfUuXlGQizET1rz1mMa54gfbFTKhqIFslMbL/q05Jgl/kNvobSERXGeB/S2f+Y
j+jFS4Lf5uxvcwiaO6Oup4iINZiLH9GRjXS8D1cqBa45+F5maJbgDmvSjAVpx5jq
wEO2qBGuh4Ibni+rIVwCtIf4aAuHeOJAJvqdKgvjXza4/+6zvVk65VnbGpJuYLte
j7BosRxzaikti21oF9yE8ivmlbSv6NkJ2ZAH2QFwCvO84dml5fYKi+I+pktKT9Ad
ZzQ6fHuFE0f/JhG0/Gb+Sqnlt/jHhbIUr2RtwdAo+7+49Wz4HjnH/ykoxxyXHMCA
wYAlVtUpygkAW8oRIhXrnxGvcnNNasLS2ZQfWQ+UPakQD8eTd/00qEaduSOkp/kq
89XMPM4C4MmsOPah6e3wZAnBpDAdcZsv1CaEaeu3CWYOROh/BZVlYHo0ORg9h3rx
xFtHdntXhPOobPb6oN8Z1GItYW0KqmAVVBOZLWOk4Yw7R+YvYbGu6I+5BxSsfgGG
dqnUHh9DRXyDGFzmOG8uA/VeNwpxPWHsHbSYVzUwOfK/A/d4mr7Zd3jnv/M4b1N/
fVaSO1DS9vY0mQMq5zsMw1L0m/dKzaMbAfgWAw3Y8KR+/5gnUsxrLyRL9ODkQXne
tVDak5G8XhBFYzl0GBrVKjMk06Ssg/q/g6Flpc8HVl323LmtXU4WsNXl36yOXKV+
LrWNppSgcuGaO8Z7E0vzg8cVqyKHsgMeN4qZctWMcGud0yqOtJo3CU07jI2VH+Dz
aGmGjqE5sXVjkp/K38BHynPA5epBAtg4QF5WUDqj2D59embATSYGkYKKVEqubFzy
CXdgAIE8TeFjK8aBQ4a+Kz8sLfgJMV048cKhV5PNEVPxNpgaDTN8q7SF5Y0wlLbN
vjOdnhi+wtOiQoQaeDYjjF+7ZZhkBvHlP2b8t5frb49mL6/VcrOJY+b8/SfgQd3X
mN+gVPZW2EuKWPkOKw9VUBonA5csIrrFKXBiU12A4982dwVmJDfaFNHDf4dfDO7f
qQW/KE9LEVbFJ/Olbgq+Y8RlCMChOYVPr7jdPjsbIEHomRMMh32lyKrb/Psd22Ax
4lfCrZi4wiBHS5QQ0KDkSNesLcDQM2jGDYap0neUxrJk73U1KxJrKD8AD6USUNsB
YAANXvRRGEEcob7rhgH3JWYcK++TpzekM5l2alEQUJcf8Ptbr5RbidnXSPEH4WS2
H3TK7AsKreq5SIH2aiEblrc7gq0l8nYQ15EW8xgKhhXLvdj4PgrPlt7eUSP0x642
CvUgWUC/rC8ozQ0zBvqGpRzQQUBb+yrGuoqqqMYaBydNO5Fg1xLKUinKhR/njrMF
6W6szECFKyWH4bbCNXa2Bj3YoEbEpOgRxSbT70mHMK3jxRJWmuad4aXye1spMVVK
FgvvXUvAvO80gHEtYMiPa96QlHd49ZBE27f7Pq9RHKIGhF2z1WMQOftiaO4Pa0v0
ZJl2aOzGRwml9JJs2CMExbXw63YhhTDc65P5Qu01vq/GcTX+jCflr5EytXQKb3g5
/mE4rZSaqf1XVwtymPvMssMdvYcZBL7Eu7HIkkk65rYN+dBvOB9tp0QQNgnwV1nK
5e1UTL1s8iK1bs2cEgjdEgtueNegUt7QRe/2veN5c9N1rKGcQpDQmBHxWEfXeZYX
yCPWEiKjirYNSp1BGC4iBTYjbU10oBJuEjp0ZmMemwK7e9G7PkpapjhMZH1gFCSU
W85n5qOB6l4w5t1b95H4+BKv2io8xoGRZjxHR5/NSUsDRvaLXOw4ND+KFQJMgHCK
WWlNYAqkhfNWYHLwgs3NSl1JMnbnfCBJhBR0IMPYjdBARh2XeSz+bbnC1PzUfyn/
Gom+j9YMh4prt7LhTazj9g69PoCG7XBZpufAWlTNXQPXAAVyk8KAfWJcx36M32Z1
dP2KjacnqIoqYVZRzM7Xe4WIG1RJZ92/sOnE8aPGBWPXGdNrWhwKp3eWxaB2jVT0
smi4LrBpisKBXUhxEfxSRQUfx+/j/yBQ9VQOCOMV/UdCK90b5iSe2Mpf3bCg2Ksz
3WqR828mYO9SpsxoxydxjD4fksdYpiBMT7JtT9PN7vcVYtV3smPhPHIBlwhxktZY
1YMVRqPomvxzdg4psB0UAYjKVghaQMFRc86+riyEURXmjmu8JMS/mUvz+ZeAQ1WH
uA3ZvxxUn/MXG0B16BECYENN8oh7wn93F4SkDT7CIZJCRcZVKgvmJc6XqCTbyA8I
M3h4Cv3qAFLV/yIaWYztBnlw/y6JxdwttW+veHngW//eRRLMQJbSnmQQItr7493t
M2CexGLsk/JqOOOuKLQwac98pXBjQe/JERuJ/jq26BHD2E8aoppj5djWrkvpLEKD
CBgekYyaaRfRxoyGrwEt2WEYgj2IVulGIFlHtWvrNKfUdpHmK7buog7hHf6Xggbj
PxnYJP8R9TK8T34XlDgrttEytEEKbX62aK9cTUW1gznLotFnSi+GF0FsVgyKvwfr
4HNzZiHtaXBaMNWOzsr/JAQGo1zTAfMvMZMK5YoD1ML8zGNIQ2iDWgUWYHM4nVKq
XiIQfIpY6RUNdjPH1HGa/2aJEDBBkD8DQ+b8znXY2Mw8oWecR/eLivN0Egg5w6Rg
87OG2CWHWZhWJ0Q4W/acXjXJXHJCiEkSEzhVeJbS+HpFOYC8MXhHxuPfotdVpJug
x3XNsGgZISLMGotbW/tUnQI7ol2JNjPli+XxPCP+5t6yVDLUSIKoYSIDO9pbe/Lf
BhgB53FHcaRe24IQFEG7lT1eJnZBGR2j0iZLDyqbGN3XFxlwaEJ4R0BMk8890T2f
dG5cWSmMcZrwttwIjXyuyKnp5O0Hf5uTIxexH0Kfu9SnysimkBTfLhQ0TWtdw7fv
FEQ6ulFwYcx/40Bk1yfA+EG8miEy1Ft2WNdGRPzDGdPe1PG0MfVI/zoZeS3JJ3vN
EP3zd1owJClrSMadX+FRglLsMLqyI8jfngU2xHxQh2gm2tEPtQg2Am/uEGmVJEwe
by9NZFbLqeDcwzUjju1o/bD8wWjfg7LakK5Qdb3PoXshqm7ld5cndd5/s+uEDXZ0
LYZvm8O/Le7qHAqPSQ+IHqLsqyHlTS2pdZ+ljSO9UbO3aOXpkoEjFh95d73Pf5pq
GSiNSOdKdK2ywbGgIZ9bi70IBaM2vIw/2BQqXw2024fGS7YhGHWyrJhIg5yRzQTA
YfYeonXeU8ovSzQ/XS1o3S5MSjAZM6mXQ6adn22USc4Tl6L+VYmKv6XHforNktWT
/TCokv06Eyg9ar40TRDQtvrtt1NYkonpH2BukiDZ2otw6GJ8V6cyMd0mzZpC6edM
wH3WxOzLOarH9kuYfFP3Ixj/L1980aA7kQE24aiDNgfSy9byssu4+98hVPN65chC
/q4d2bG0N8GnDKY0D1h26RDjccOKHmKgiHhje9KdqSXnnRGpHmyRiwRGxuAg8053
8ka2My9po2MO668jx2fvQf6DN9F06GMV0koe4QQJhEyH9SLCk6X+AQUYRcZNgGZ+
dtHeu54AHvcwpvCNuQHsY3zKfIzRH/HPZMgYxtkeCJ/WiHkuXNRSBFeP/pKY0bxO
/m6xt3/8Ak2GgdQruYS5O0QVL4TZzlHLAk0wAiRmzSbhgmJABMUj+pxZWlGDzMW/
2H6v5eVOOT9yNj6zWD5WA9W0ry+xv0rO+CTKTzXsghIZLd/jD7oJZOCsYmDBQsk+
A8IpL6RoMbwym8x6wNncqf0D9RDHUhDsg/Ug3HrAr/nNFv8rTOfMqzqb/tMTFf9x
kVeGj3cRn2BtMY7uuquvAc7wim/LBaSvcOIhkgRjYVYnQxDQhdfebQlB2nj3Vmt5
zAPYVascwZqkGC11E7jQseamnhrcf9w29JODs2vfsgiSGLytR/c/ZYQqx1D8h6Kp
4QgsWJVi/uq6TbNwwCz1W4zT/oqukHii5tX9MTcLVmQBMy2M6S8EdEEbsSKJ09ba
HdHwmMGCYO1FmOHWmAvtWWSOmjBz16kj66Zo3TRN6HwbdpJqezSM0FGSrfe6rIdN
8s7zXk0qgDyewnPPtESJ8f6hS9jt8WSCKMLSR3os7jTR3gdKo4bawIAYjAY7KwIH
EUsouXh7dQFu216K7gfYyBpo8m0cLW/9Wyz3ZQvr7B0ToMLLtqDelSUa5+Ezg6S4
6PdOxo6YUJ0zpd5CVka8QT9V222wn6wpqKcRBAKHxtQmbXpfFY7Qj+BI01X5rIyQ
5aAHo3p0nKhF4HFJbQ1A2Vyov0WS8Eb6kZbm6EHxt45mBYkTJsJrVK0TTtkZiD6X
Fnu02RZNylPA7VWeMxsKld6stkRHpI4RP6SJyB/rVdc0tpU4g7FTqPQCS3//b5Bh
FSuHoxk7g21QG+HvNe9YgS6wHhfbTKZSqo2Pr+h/ArR3LmcDhTEcCvOd1lCJkdC+
zQqDaYm4FhlVDMP0azwrCK1vp9FNOZFgD/5yxrI8OYbJfmWixu3pxnTK+6cOhtfd
mNrQXfSTi0vLmPcUTgtkLVZA3/h8+VsUPCc3JDZUU0YE7WXs8ptKTqJOBMus0QTt
IAQtHxCQD6822ERj7U0hOZQtnDyjw6KyurBqCiVSQ6EVDLqYNU8p0FVptC0P/TfA
2KkNG4kwSK5PYB+JPTj9UzOTGRbmkNsZF6rBkZVJTUfVGWqP1OkFhCUS/72eGTNO
VgB8z+8YmQZXCvUyPa+F1OIOnh2WtuawBkbKZmvGgevmMr4A5O5pNWIwzTNUKQZ8
m2a57DDKMoszmxwzYotQ+XLq/V1xi1HrZhDPXUk2DfPGIY5+mWBBYWZqVy/ReN8w
QdoS9h9OdYadCnPDZyG+FNZ5y5l9xd1g1GeD6B6sN7zNOoitGQ45aFCMWL0muHjf
htcW3ISFNO6s/9uRQesdBCoRbxxKYKzSfKD0VHigvYgGE1uXuHNYj7PU1KOev0VG
0C99fhtxSRMui6I17szbvJhV6XWUYlfNXdHlAvlnXisDPcKgr6G2KG6kua9Ss8hj
kKZXFJy7YXkGqfd2CJ2TkH9R81qIXQBTSxmdqewONyAmkdc3LAbm/sLKPizbdJbO
jBFCVHtls7K4fftsDzz5zPLtOz8FFkDiTPY8Vy5mXjVFl1BxgYq9zAeioHOuWkc5
h0Kl5aBdAGZlKxPLxp/wRPEt6AXq3ZDDKdkOBd+ppucTcNz1iLhoUGfhiksYxu8N
k3UnJNzTVmxSaa8XtK52hz4+JCHi/DycEEn+QoGaQ1MOxcExZ5YOc32crnl89QrX
0WfojLxg03nAQihcpqK457GrdHDX+EEGCKx9L6ODyxHsOjKuwv6S7NNjiSP0xCIK
G4YbDsxJ9mD7QsxFHhwk56l4hkShZAnw9TFI1NZxu/QJdODjFluxx9DW/KuM3B5V
AkZMNe6kfJjFh9HqTxd14CqK5QN0sVJKB1EUeUDIQZCAdcigA/tmFxyVOGg0qzyA
Mz7JtPAX6jKFbeIGUS9tz3lK+T1JbaG6Ia6uolovQ2sEq/duVfsZT95iSglMQiRY
TgQaZhFDLpZb2B18nFjHqu+mo0cSsqb847ngXcmaYArpGCYp0VRNDKNEvnl5Qy1A
fFrLJf+LOmpx6jG1D+GRQ8dwOwqObwIPiYMiiOSkqtwxGZ6brfZ0CsYU6kkuF63g
YnpaZJ81E44x5swirQfk2NgIfaZ+Hy5J7WGbOTSn+JDpy5M+AbM3wApa0uLdWt1G
vgZZX+/yCawTMwlwzQgLigR/AW4yBFi5xINBWe5MdCTzGD7ukH3h7/oRXcc6q2fV
Oa+LRwmFJmNnGdM5by+64bRV66I2taJ/PxTRwoxwNul5YDUu3thbBFghUA9WoBdm
1ygdVEnE2ltjyaWh13RK0yvNLbgvnX67WSvw1pvIcd+YvopHtcXUB8cWpQjCxGvo
ANQ3eVpoj9ldIxdR6bwNNOjZLrlngLwaCfbVsYY5M3Wx4UcRT7nnyyZQfBjPpNbS
iuAawcLnUUo3+tcPLspNdg7tNBQY0GhBSVqYFjzpUkbHBR4SM2kTrSDpfK+3EMIM
6+x0OPCo5EOcZNfwTXZVOFfD1c22AWpZh8VJ+L14NObNLyVGRNyvAZjlFuoqDNyZ
oZyxoLgOpFV8qBqhMFTAecMvxufl33LApllyaZp7j659zucatIEF3gyRAuj/tpYJ
dgN79MfuBgcEf+DpPFQmPmhh3HxvFkhs9vuAU7SxBkFibO7+S+s2PrXOQCH1i9xA
bej5CL3bYXN9qK8MH2eU88qKCKyQ82mj15oRoBVyHrBf/Q2/7PvRjdaIntNJkKoI
qf2qaOJFSv05jXzmCma0RbfKU7h3/S0FbhTxJTpFMWStU4ExE+8L83aPEnkP9IJS
JG1Ky86PKVsq2oNzYbwDd+g8qBjqoXQ1rb99K0Hh03gc3nQyFWOUXOuzs2rdndGj
tXWWA/aI0QjyL3PGeOJ8uNa5Z9wXHieLROMzrevam3b7b6mQLWuQxlMhp/U9fbD5
3X76iOeWmIzrAthGA/UmNUBYIABYfI+KR0gxOg6+woPz9OXXWPo9mO/JSRz5xRBo
g+L3Mfo6BPT5Ji1LJKjR5s8X+aU4jlJBUa7dnS7Kfs9Aje82Ks0P3xb9stUFm5v+
yVUOFgdQYsafQG+q27gXQBx0J3AeMQk2LW5VDTJbK92/v2fIkXnRpfHCe0PJ1aPJ
29IfAWuKeeK+diexYktpuE0m0UJWVl3auMyTYwYNU+jtH2gzBH+eXM3BCqpg72JC
LV+XGycRF3A+CV6xNaERqOjMkYMLFT8AQUiK44us/NlRFA2dSmB8xFCqJ3xEsSZQ
C7b5Tk4jjwnimxIhpipq0bz5H25vuvGb04Sz3gqYVx0y9hUHO398Xh5ta/s2Xmbb
r7HtXwZgNv2C93UCW/xk+L8WL772VQNWMfZBMs9pJwwkY7o2p7D8fNJdgQCMSXZ3
630vPJ/Db1IipduRMlG7j45BHeBnmBXj6E7mq1pOD6Bn+a8VSnfHsyaZbf80k7r6
LSEfi/R+0jtvRpUzSMvp4dzkzbFdjH3Mv/5U57sGfpKSI/csauFrQaijmRjFCM4y
nWrRFiG3EZcMj+hnDu87RQXk4FKQWiK9xXuq4YnHojR/zZZxDiObukAYIl79dbE6
IaUBmVZ2UmzMLBGVLIQtOPFPVaVcji4DGQx5/PuyW25Dl0aVr0VuQwqCFZeHu/as
WvsZsoieBMTgo5eIhaeVW6z/ACxoHtKcOiABLUGMQhCbTWlBotjiKWeRL4KIIBkI
uhehglwe6e9aLSNfchPuuG8T//EiW4d39c6PvsDNi0oaGhjhb4rzdd73368H7RJA
HsjF/aT3KKoCiLazSgFWS8Ugyl94Ma1S9dJD/WqSdiSRxW294EwawthS7MccAEfq
I1GehK/3AD5LoPKnJ5QiJ1K3gIdGhu8h/6lpk3h9B98e9ozhWtz8gYGAtBrfJH4N
L1hioy65KRWPZkCLVykX5WSzVMP4nocad7GW8GEAFZlsOfe781jCNeD8kWl1jmG8
MFlD/FfMfSeNJGOQBzRotKIPZOxApbrdmmkhN+ejopHaOqGu1BXIIB7ekSuYzgjW
/UugDsCFWpYJ39mnBAvNdQHSZD9+MmI3M7idhRzFIZtt879DKO4z7T3O+M/xO6KS
3iCo24axXgEwScf2XKAbyXDurtr3z18nRciqpjvmvxcQscr37YhamYg9YH9d7zGX
OFE+pRwsgivGxCnUfwinl8FkZuVJhMwh5rFM0FWDYA6pa3gi9kdVnONBLdQ9SRBd
G1/fxf73pMmp6lXE3E4OPW+f0+HAWAD0jWXyrKGHqIfvt5l9XNgJ2DJhTphPaAu8
l8tA1DEg+l/fuXFwsM06YoYXv4Kgc7Slnvepl3hYqBYEr5vczqq0VMrDs3jUzscK
D7sq3Pow+Cv+cqiaOWXU41CiAghYgXaJEKbeb80GyQwmcpSyqlC50hWmHD+FcSI2
9KbN/OntE4jyVTRjL+I4qUyax24riGfzhJygvqOnaZE0PoVp6HvwDvOoFlWbNpO0
5FF4m9yafushdXM+Ez4TMucCZlRJdE5zP9h3uNKoZjf/S/4NCXOSdpGP6x7dduNI
3/9xfGanvJtXsgRi27BEqYtnc2wPiu7If9XYACEyQQLVLyAMT7qfk5to5dUiQmgw
uYDcoP63gx9yONEFioIcxzKJpQGUPZFyxQTatvAMCXQG1yqpXik1+BDbVFIgfK55
Ql+X6+tDxTmEWYEonkDHdzfZ2uR/jK843j+MU/H0jNJ1G6cjox7JXYKTLC1cEOe9
gvK+jt+vcK8q0kNob2JUmMMgbZ0E6Hw3Q5gYYICud0E0Q9NqEpJYOhJkobVrHogM
xR7aWv2vJg15s+IfOmii3401FoDTwoXyGJ03fxs0hIcvFFA+RlqAumYe0nu0isev
eAWSg7xEUgAbN/y4qTnTg2bciakPLwZiBkZUzTj2VuKMWU1YXqvUDn54iEvodaT1
S4OkZyyYKnwNZl64EeuNHSND8rzLPkbkvdVKihfKNVitsctfJyDk7WjM+QFcyGjE
6SAXfb1sZNOAL5uBDUQAzSzUko6DsQYDRhUIOh6u5J0NZXIAR3rlOJYKgdGNEoUl
weoJMZ1Ge8ZVCChq7FyQspwduo9LF6H9gpqzqTruGNTYtaYR1mFbzHG6P2dzlWz5
97Xj9Gle6DIzDgaupbfR1AxNUlMVaDZcQpXDtUHSOeu+ZjRvm5Uxu8R0MEGi1efF
1hWGeU/F9/q0lKKCDUU0tVazLyIH9moKkxb+eMhLn7lqKdyTQR7KiwONab3bKsWS
21UIGH0BnNbCL7ILXC1ITZAiojjbeL9fKpI+37X/Fih/B4yIRRzNuihFk0DpLgMu
a81K7opwKvtG1vwdp95TPedfv/PwplsCmoECyeKDSLD/7URybfNr2NqlcZTLiSvi
dUtn3gWcbK5pGXjpRL6J/OJfe/7z7AkpzOYZmgrZvbVU8CFLAsiJaPkMHdtrvOOG
EjPIgyln+hgM9YbcSLEIHi5PxvdmmxpD6H03/E8Rz+CZQRnZLwQ0g7j7kws6gQdV
CsbRfgyNCBnF0ToFPDZy9mS6pTVLCL7u9yM2H+wLq77/n0tPndgwiZLfoFla746F
zyHootREPC67vuSx/g9q5qwdaLVjtuDxFPQBD3ADE7Ts0VRq/vaZJVobqaaO4Q/j
Cucg6olHL5hnJUd9acbdOnZsDo6H+AwezeFRniYUilUxjcAnYMOs7HnnhYqjf1P2
HrDqfk0KAtgd9FR+VT+Vfiyf8zk0MZqgLkFJdq1McqS0xtPOrgaDRtw04FKowE/k
Z0f0AFhSexmj1b1w2BIzxXK03yDF13yHTGTx9hna+iSzi8hZDY9msM7LWEVy9Lse
Wsajm+Lt3eHFm9CKBiHFkeqX2xoQ+EdKCNPRPHcOn3HlT2n3Vw13wKc8tSC8xm1d
plwY9NGcqr04D8jbUPNzdjnuxQZohvGXjGT5YVKtwsj1h2+AYzVvr8Gjr3M1+/Cv
Zs+6xcR/7sJeiA6Mr8Ud0HKlstk+sQIOeCu/oV+wzf2FmAXfvMdYSgt8Dp/1Veur
Cu0KrftzfHvgW7GoRvM8bXU1WV/iKpXOJ+v35L2hEqOgRFKIoqHzk6VNflhw9X0A
AwcVR+8PZu5FnOhmKkJQfH5QnNF2g+1c4kn1L7KNPqnRRVAppyCzYobIzs2taGDn
uOVN1Z6FJL/xOnmywSuGsipr3crcs+bvsxuY5qj3Ah5GLaOCwrba4LdjYpqlUL0B
jSiPv3KjxDRo8b4ZyW1Jb5GmokGsXb9A/OlvWRvGhaeJa5VmC7AG7gXOsTxtUMOh
cyfBs+YJkrgoYTOqFgBnaYTZLUcJggNBjV92tVE6OQv3wytdciJ5Se8iIw3NLag9
67UUHVVC44Rcdga3Kj48KLO+joAAiQIFAfRzKqDbtNlWgKEvMIIMpd2fY+Hu5sDp
Y4zP6hc0YbWlHz9VgVmcBtGFa4yo/KrCNFcCaIToIPRqQT60jqOiKjUIBmx6rPB6
uaaoUtMF486ZjitaQv/NVHumTjinAO3TByKeyyFvTNV4Uezd7qY6NfFI1au2qkTf
3HQSeDtcRqfx3iW4pCcWZmmGRe5UFwTyS5PmNeRTS0b4idiPYuIySQI1W2XjNmSV
fKSc3JWgJt6oRICvWisRMwmmUD3vTbb6NGbF4UJhZM0GD8Ayv2S7ZRRjoTQhvyGX
U+d7e7OHcm8VU2KwEZakawrn/rQB7u5lxMKA27IREsIK1gIBqohMRRftR23WlFmS
hid79nlGMr//dHyRLgI+nxIBUuuaYQvHiA9dHuONuXEyd04yKY5CYCWJX8eC8Drh
0yqQbu9A1JDlVJV/ch8ocros+Twl+8uAfNSVXlDjExBmu+hJfIg2Bwu3eAZhre1e
RZc/lV/m/23FSniRaEa6CUytZlyVJwUNQrjAz4ZDLTaSR71UXKHsgmYILambecCv
GYCTDmdJZ/UBZXKUETpZOmtLA16IM6gSZ/uWIyiIv6qCrW8Y2MdxJYwhDr8CL0LM
J1ZVvvhbaLlBaKtwWv6nuZLmNOmdPeN6dFy/4osUnIX2Dv18SQP8PPAOSABYFRmF
6q5ly0cS2TIvsuYp3yaii+Gxu/19cyhrX0HupBUs9ZAQxCzI2MN8b5/RoeXA/Jdg
SK7ihb2ZFGrrAfHhf2IiNHmS7No0rMPpHHR0hldpnCyGd06ml6dpg4/PR4QNLJ+C
gbxMHE29uvlINkGlxrMF23ZTYZP+8zrmbLnveDBnUb6oBEP+c+E3SblpOjChF/vm
CMUcjkpXYqZsFgR6tAuYyIM3NqCyD4fx2jY1kDDI6N5cSj5FGFu3JqDKJMhbyDEV
aR0kg1z6tC3ACLWrLJXKyYTCsjnYeNKEIH9dCuMw4ml9iJfnZKjyofIhs6mgob4a
p1MfZpfk4yeB9pcG8gIJbLUWoDl2QE/U7GrcWBHGwTCAugXyjLDXvXfcz+s1PyT/
4Bgi7x3AMKBbMLqQGpSyIpCgTCF62bhDebh7bxBTSTbvxPKx6wdJl2gtULvaJC8o
B1AeR8ohITiv1uoH5CYOopcYKY/eUMulFTNcLs4etXLH62P90MHlMmosGNm2VkSA
fQ6yj4tqCyBDtaCfzdg3lROjwFw2lqeFVrGZjj+appKY7dsj0xz/wSzVD6du7yqX
1jlulpp1iOuqHaJ1bRFqLI3PmdkBfIXiz2Yal/43I10lPJTv/f6z0QE8jnr5fZ6p
Vfwi+P512B6NhtJrl4/+OO2rOqmkkM6PdSBE77C+H5PDzhRlE8o3X3HrQsE83rlU
iickYNM83PNOu1KCN5Hh/8uc/AlmfFRfX0HrlsBBqub9FDwNW02pTTwT/cgBHaD0
7VPsdar0Mb4jIBTK/FtwtqM22swLA9ru03ozyKX3hFrI7jAPws4VzgnIMTGJfPpR
ZxUiHH/f7LggN+DEnydUL+J1C5t7Bbr6EauyajtNsKBQ0KmCWqFS70e0L7/B15uO
SPPDg6k8WesMj7TrmADGHOc35chxXpQmUXqCDbcuxm9RMZrlw063lq8GBFtrJA1B
C9r9KKt24VkTadftDXzPx038kFRtwap+5mAf4x+qU3LdSwHTwGw4sL4h8o28ZMaC
K1fQJRVOKJGNXc6iFwUTB3UtbOj/v9qFTRuAZgxa+5cPpKqMBQWyl7LNmR+6Uzq9
iZSqVQ5uMzYt17JvCt3yPBa6cPaziTurNU1VSX0O4JeStx7VNbLyt+Z+rFCqotIj
xXmVXqTAd/itwmIik4SFXFI+aENNSMIyT7/H3QZAusOswYUDVsjo6+GdxsKDQsf8
3Ztenado9cn+1aFXxA6fQSVefkCNO1J8Kk5ov2ONH6m1eUDuICjiFwRh+HZ1Enf7
pKltPHzCcB9rfJ6WarTYnMm4oReMy5yiC05/5LoN0Js87J7Y4tyUpiIXXUyo0Sdx
beT6IdB/a0tGXgV9jvoz3+dfXBwE74KhXHfqLRvb6JA3r4k0STonMUbyEBX5QVF4
jzdd0DC3XRMxjkBaQhlm/9cchY48lJwYWkqLGKyZg8QEx3OhbuDeMHicmp43Ajed
NSmhTPW5hn5yjuJtSenq4YYAmn+iS/tCSKTz3MvDUFuBejD3D25BANl7M1NRZ0eN
oqV32gVs8xhuloiznjbW7CjnoGJUsaQTewwCCVE7n1Vpd8K5jMu36FhsbqkP6H/K
TayZdkATYxXdlLJx+fDvbWJEexV+ztC1EA2gL7eiHXs06laQp+pI6rtqWpttq/v5
66OOTF8bVgDAmqGCPl2MceVdGOQevSL9FCQWcx98VDyAj7tjboZAKLaD1gBKpE8h
ahkzosqz3lS0IUJYXhQX0mmH8cYTkCOk0M9zeCruZUfKgITrSIJPHiAmJ/qAb2Yo
7u528pLxLPiAdEGoxvKR4OiocBsyOitILKqd5+Ion5D504vY2uD+Iptn5VJ6nW6R
GUeNBnzLkMyOD3B0PxavAGhwJW2yIocO1n8SlL7L4NW5wM6iup2/5Ge8Hfmiuz2D
yfiAlXrxty/RsblxmOBLGIZgrmXh6PmXi8rehy2Ntl5wbQmRNKxTHWuzhl3AxOaR
MDxoibJIbuqIZMHpr8xqk3G2IK5I79m12HJH3SUQxLIYvt/LcWJykPGt5ebdW0nh
YsdLFnKOQ5gJRSYu9x9P+nFrV776ciwELEUn+tiGNdUsoIoJYTC9XF8thwNHfJoe
D1MX1r7cYp5euJtJh1XWviZ9AF2S0SNNQaGCyj4702iwH7g6fcBd6aO4ZxnSapNZ
ea2JvFbf0jRV1LQIe6tn62jKBBNKKTT1zyRcxc+cxiKaKEid1fyeEFjFdhwWxC7o
FPdlrqz6p6aHdIVfZskFNn/Cj9jYa+98ijOi1RrHXLvjqot/Ca/5i6cv6yioJpxX
aAo2y6Q2XVJ+i98wqUi245zVJb32xuqyjZoZapUPBjZOQLq0mdtFN8LIt/cqpex0
H5PcAm+oWnQTEdI40bVUQ2oXUIjS0HuBX2XvmYx6IXjNoXTNb5cYbl8/wU8M3sk4
0cKhKiIhrmdn0G2lnXcOy2vKGc5eMkCbsMDZp1BImg5ms+batRjxFnmkmT+iOaHq
3JA3kHCsw3cI6huMPRMe12+WnRkaILrvPNMcIipFcGwIa5gIAJNGzAbv70+v69s7
I75EsaemItT9SSMlHEOQxltlePOO22JZH7t6WP7Kv33eWjVDitynq4IKWCuNEx9u
6hJW7+h+GyEb2LmRIsp+Mtu00LREidHebMk7pm0p0oaUDMDBYrBy1HZibRBNtPGv
2r6EFv17U01uwf/uknH6eVfWCPVXD/W31L7hK/QdWH8JJOzgmomTzCGgKSuP7Uxn
uWoAj+ChKVmNpG8MzOC5C/V7cz/Z6yY6E8tnYQSWOrv6vkPcLz9DCMAGsho71/14
rv2HPzAm77uW7iQlteCkdpLtGSDhuwo/yr/82HnMZFd1+vgVOUlWBcX1Wl0kwGli
qEfK6nF+Nu2oOgSZIxt8BR65b2wSHkGqzJ8s2jr0nnTY6iME+5wAuoAZyMPTXlZI
NznpyqXx3Y4dDZdHSaJBeMaQhXf4tvNsL/su7AvRAFwO4PX26qGqzUiXT/RjVEJ9
ZFBRB17JHTfbXFEzpVar+qAXh/JBdTYD+8bUzQ3GMwrtMvX75p/SP60IXEm9Z4qO
4IEDcHdfcQ5WEB1eSOaM0D3ZicQ2Ryrbxp1d3BXH9+NncEmlxJRGAjZh+1JmcFKH
+T4Ym73ddwn6x2QaE4LcIP8kngir/Hf0D6MZTc8tUxCPRjj0GpzUPffbh3aLArha
bOWaYSsDD06YUDQfTuKjPltEHcMxp2zkrhf5WPOkuZA+MyLrkhl5NioeadY+AGaS
kKQRVij8ZCr2U5PtXyXEBEaCjtcLRPZIiZXtcKE4v6u5QkzMw5cvxK1CkFwOaZph
tc79tByq7546ecodm2bccIrPqr4jjmF18TL1PvXnY5mjdTsG8o2+/3bv+5ARyyfh
VM12uRdjMQw9fEWWVlApAXt7Pdw1PLHmuL2HYAgAbYGUCGs/ZPZAbZlF4r2sXkX9
HwDN7IwXzr4rh3Y7w9DdWjy2kVPjivbftGnk91W7Qik9YdGdNk8DmP7eAPvv7O2x
oXQrOdpp7YfkNndaxAXdie7OyyFq6m/x5keYIqk6ijORuCc/f9ouzRzWLZkzWA7X
ZgQQuboG0WRQNfPzBYKwDiYtHRzUj7Y0Gr+l0lk05nqu+Lku1CM9e3HHdaVlvKpm
0s2yP2tTZhTeGmUpi28yhrAa4wBX+Tl/nBVFepx53vj8XvptmypDNa9UtAWyapCW
JcxGsNnl0W3Vc+qBfPPRaV/2VLGozAiOtVhVCyz1iehoqtp1nbikZ52IbH5Kb6X/
zYd6l2h7YNpeRJgwgf5pluBa86NeiWUt/nIsaISUBQB6QgsZP9scomEov78oDHdp
w2WWHIn+LqlFgDavmOrFpU1ixItYfMOn6T9kA1DcAAS+a1g34DO3IgZye1eJwuQ4
/D6IOscCVirELnLy4VzfI4LwmRqfDs3XfXzfzOmBSkvltEjdoK8zEg4+BpkgDUDe
Icu9JpAmheeljPkn4t5HMfeMFz6jtK85gRHapLR6Ua6iU4xEAcWIn/u3q9Gwg5Gw
lnYOMALrZawWxZpc5rzDIN9EB8EnJuXaBN9Stj+0AhtueeeOSzd8ZvYjDaS7yM3g
K7i6lPZhrX9pI8ejh1iHjCdyY0LkvQgBTmvPxhz7Vf/sMWBvQzzeYFlcER9ioKf2
4bfP64Kvapo60yrG9t4KkoWMWtK5BsaTbwiNqM+i65HBofd4Bc25O9SJ1F22KZ/O
XTyDkW3+nhKY8H1WyPeMhhUnV01okODC15mmipoVofa5K4LKVOaR8+Yymon7xRmT
yeRK6qpUiT8AprX2Vbj5dwjgxH1PCYxfGz7Vxa/sRyBmTSF6IlzMssvVmg+9wPe2
9eHcJJrB9A487xUClJtHeBaWU7RqbaS0n80zchlEXy8OjWTrV0EjwWIfDsKlg60F
OrdufvZyyXnO9Zz1/I+MIn1ZuXTGpQ8zKtGRF9BiGDem0WZ2wttUJPsGsyoPd01d
N1uv/ufgx6930DTKDjNIA/Xu+fIPGcNVr1K18yrTqSG6tgcPnPGNfaJZn3wxs/wr
G5+c8Yige2dsrdz3RMDLafumEC/2QkD2UiIsxKNtzO4gMxztJCtkcWxGQXqTgcuC
fHmwqkqcH93X/9KyMWatOGwJXZtHdkiKXBOi4Xtyiz+EAg6BXycjyfMsHFL/osNa
nlZ6yZJQJcazPsKzaAchJEROBNVf+SIHX0Eq8vhzQl6g2rvCIYUeNz6CGODzMH23
8wQKq/ykNE912jK6rkvmGhojxdY8x7UnxRYsoAX9b//jQHLzsufcKWUNCbp50fcd
pTWzLO+c0ln+BxAt4TOnQijPm9TEj2hMgrOV5hJdzrqX62fCVkCA/k2j/yiW1PKz
ie0Jul+YCAn4Q7L2D18uhmp9a//jbT/w+/RKqGksKC3zBUUvYvC02HwFXzjnQxMG
/AWbUrB3ZOd4iMwtphprnmbdYuzDkx2ma2AISnxglvLrZDUd+HQ7oXngIY6WML1o
t+K2LIYr/Lfpv0EdvMzVrJppfNwSlZ4Itjr3yRc6b07gSjQX4JNZJNQeCCQ1TKs+
hxI4Z7cvg0lvxFwz2xV4x6ha/Bd4Ket628bDrvDPbSJtD4em23QmiVg/dl3tUNvM
ADpop7l7Z1CrEbUcpBmhOF6SxgaJDToZx9KFVtXtD4UlsVLaLJ8nVSGfxZE8JPS4
69/3XTfe+80EGPeOH/yAaxXqJLTF7eOoEv+kZ6D7sbaArmK3325CgCQCu8HrLc9S
VDsQcfrV1oZNJtpLzMfFoThiUov0bqR/wX7McWoUPqt7rOaDZsSzHesgkIQhLzAV
1CXwp2rKjlsT8i+tYKq2CFlyQkNqm2pqiFZ5FCRVeNBggWAXM+KjVjWkqjrCgWL2
YwEkHQ2VYZ1Sgq/Kj6IE3e+CWdWlS+XZbWL6e0oEOVl3UZjRQ3YWROQxFMBnJ7vh
8yXASKb7GmXrslAbgxaZe5WMUgt4G14REw2IYjFO0wtd3Qac6Fe802klQXzr6Chc
Y+EdubwoHJH9EJUMgHTE/fLz+YoguwofEFcbBjj/ugVy0M7NxtZlSwD9sUMD+gks
CwzlCCwIgEsImQ3YOrs7qSawHKbjN4gwWCV77rue0O0TtdKtesY8ymExn/RWpG8X
1UK46TqCD6ETz6guYvW3ky9ltPOZiOHcmjYjKy1LWpEMh10/jU7auWqZznoW8zpG
8/QfOWwQfy6t49inxn7uDtCXYVNxOIsbi90J+oOl3aIV+Uk/lMO/ID+DAiO5AgXL
ykANPnHeJvHYd/3PW8DU53nBcfQDHAKOWQWThp76hPgvn71kTSTKSyBnQ4cGgNF8
d3d1bZYkK+hAzdgy43eQHZ+BP6ml561fOyYKJs8uQL6rb1DMqZqqetqGshB8BND1
tHurM95K3KcyoGlFzMjzKtMF73ayLx6OZycXYIrlJnLgTWRCWk1pVjauN+WsGIPF
WL+eQdnO+omaxoAgLjWx4FYsWZG/57pR6iBhj0Jm2wOdk0kleSypq6SuMfaprpcV
wAAUTp0e2HXfkyEnyOSYZPlugp5I/Svfm+S8OnfeBARqvTDv78UQIaaqBeyIKWiF
DL2QZV4IAvJVxphZTT8ogEV8cuk/kGeOm2Lg0T2h9CfHrtMOnldhPi5UpWor8RXI
+ph/uVZWBl+cdap3OqgDMxxz7SV8LITn7GVUqqNJwLOwqPnqNp/cpr1pLi/+AkmF
IiznWA/fBfSqu1Mm89WjYCS+6yM9o87F5ZDLlo6iVD0fF8XwQUVbacVA27H/d4t5
7uqytqErpr4rSsRNrYcv0ssteMnA1fmUDbvW5Evz6fMypkWx8OGaPu8lgXnSjGk5
kdS73q6SMpJ2YhTVUfUDOBVPAnlUdFHpFnxbAkk0eDn2NQRXZ52W90BAYrxsNyyv
Yx8497CT8jp1pmdcFr79MrfVG93Itov536+deq/H1gIROdX3A1HCD8zu0eAT2lbl
OkUzIDwfzzIxWo4hhp+0kW/o8ndFBG2f4YJ2fe5diMMxwBbWAJKmacB0Aj/X7lxH
0F9ZQpiYMarEbMnc1MDCiG8TMaG1qCd23OQ0MN7A5S/eu2M/HPJSuLiWUkoB3Yyl
aBG8PRRtghE7YMgAVbS/eJuue1BBK1SYaJDWRiwlwlAakxrVxDFx9viDe9mLJt/l
6SGH25fFQZLNUVBtlUcpDSkF0JfyTGhFOhCbD2hH5Gf8G19MuqovJJ2OPEeKQFvd
VoBYv4GDK+JN7oHSpixRLNYZZqdBcuDr77tXuLq43bvxNbw08xcbCGCi9VNKHzpZ
IC7hCaPD0Nrg/uMFlMJwBSgjQbKoZ8nkNDIWYBKv+JnQMsTR5Zq53oEK4ccaa7mn
2nzDdqu8YoTPTyNZaGW3+1IBhSkb4IxfdScojJSOIYlfr8BjMaqT9fgu+ffgFDzt
cXrwNAYq7cmDNVhpwZ8+2QbEyguebM6VZBPIbOLWPC/ySQJwmYkw3eWI76QfpA8P
TG7G4ZSJ5+VD6ypx4miThOm2C0pr2wa6jdYkdRTB6o+rppG9oJg4/M6brthww4Xu
GWSb/wa2+e0s2LTpZyiYIDuG22VsXUzhQ8ys1riy6icKh5kzvF9eLswWarSzrGfU
Edm38lvs6C1xWYKmTiOw1AhHp208wM9ztyqHCfgqoJ+g4HcS7Bqgh7NRqv9i8WaF
RUAtFXbB30kPEEo939ORLovMLSQkS0y8fPb4vpsaTP8vEJpdS+RSbx/PNBvm6Bl/
hJfyB2+CHSncnK4esvzEEhagZf4Pw4/XwXELaEv+8g7eucMiXnc7BP/XWOXP8Ibs
OOD1OigEhwbQvV4pGoDNOmnAULsR7LQ4ssR0rekivDMkzFQoK2JJncsVqQsfYvct
ucHcKgjTAPDzBEl4gCPBTUAu3gV8HiBb4HwzTlCtHhU5PnMdGDz0VzhDd7Xsk4tL
oKXIkCrFn4F0n9v2sUdRNV9hNtBq5uL4tO0cUOCTKBX+msa1RBVRYwKjqqHATSwh
oYLEZucTScyigZmqwQpyfapAjQJqpjuURkrZyGSNXwdKeYzbdD5NjXIGmabjjtdu
VhyQswhp1DMIG1igOpq0vuX1LoEHWK3ZncXHSOyX7ci5QRqeb3WAGSH+HsxXIKsk
Js5hN/zycOhDOzCQTGRf7vSV1cF/jWHb0qK6esiTgZ1zEdKNFLC7/6/kivlsyr3Q
GHsK688DYAvYtXTIUBUaoPcLoJZ4wnXGucwDvfY6HVR8F0olynCinf2L5DCyMvbC
rVYA5ZBJFna7KSxZVwPCNTiQ5lnkEMfXgi/WycWdHojhHuBeuJyyAeC8X9o6uxYG
bElCiXXbxt29mLK36UlQRJkHH3CB6OM7EV3NS4IFKeSVvKc+Zis4roMt43hJeWT+
bzDHoc3dlQJzuHGi+pE6TjQ3exeSTh2Pqb6I3tHtH2iFb6B0rS2RmP/e67jK4TSM
YRepFVlWDMHFJir+sirJYjUitwknzJtKLsfOb4do0YJDMBlKxxhmuC9bK8YByv1r
auFq3HDDT64RrOYBIyEph0ybCBKVYWQ/7i+TBHSo0JV3esChRe3VpZ/wvdrcE2EW
BuevJSWrLSBRNclxZ9bSZBOszQnqe1DtaHeceQZkOR4nyAllKAxFyFRPqX/IPpbn
hh70OX7jf9VetF9K+fCYDAP48ZgCh8Qb4SP/0qYGG/uU7xpneCcxyBuZF2Hl+RJw
IupExb0hG6f+BOY5qYkCPK4pz9nm5XExQt4ORvbfh1swVhDzBaCD6DyLxHgE18X/
a4WDrbBd6o99u1SBOQ/BaBrB4olekDuHnV/WHCBaesA1xz0rhsWU6MLbjvWvpZrw
0SxTkdc99yA2Y4AD0pHShj83r28oVm3CkHUiwT0GWeJWhMKVLtILiJ4VyIlFgpL+
emjRMqWdJl9R2oVxHw9EcvxrYZ6U6sinWwX9nNDNjAdpO1I29CoQYh0wFg7VmAjH
JYdu6r5bE+irGZDjmFpBmlIDuemZQqR6ycW+ng6pkbekPElL6NYvCGg+bvbJ0yuO
lH5s/N3Wn1xhqCWkbrC1mNEls4Ka+hORtt1bicRcr+mfr2vIP1T5OqpKRdCXe+Pa
bMFrK/LuObKqcQB2uqH2g1XI8bSU9gDtDgJTOqUvexaM2aIYnsudho9c7VXushXC
1x+4ytxHk4S+9T1Ke+rJlUkokUz1k8ojzuCtmDund+4/n/Zx/s0NigXEV9o9Wsbc
1Kk/bVDa6QRXPy9b7wEC8z+mxn97oLGU58I2HfNOJD3mOjtxj1cWQBO5nEEyEIka
JF5jLoOgLX3Ffx2f9YFG5aDnO/PcbMowf1C7K+1KzeC2SXJoFQMAfse6iFcgcEoy
/QLC0DPaXXFd5CKMEwMcZwM1MG4wS9rwEIrPeD2Nho/xxAjumEfmRqd9d133xvxA
klYCUHJpjIb5yVmC1ClHCVZY0wzwqzj9yy/iWgEuBdWpDqDkBE8EIXT28KX6jS4A
Wasw/At9uf1ocSdCMlwGdTBnxTkojd3j+Fms0iJnLaXF+8214TJ7+2OUN76/gmZA
SUYkEZpS3HUHZQWvsWFC38MAVjAe/w/GjtAgc9mfIVx0XayaIYc9ZKGXzFDYEMAA
eX7imxzbJyKXNCGVltWLDbXmxwIeoFIZXEcESwkCqY/QcV1vzg6seVulOWalwkpd
OiF3hWNOIYkwk6GGupN8IBCV3vTU/k6qiuLRBHZPqY2dglfLLnf73fzfjsKkDlp9
KN1zyo8uCTbCrAThBeDTDz0LNuQRd421k7PMfyegVVZiDXenx79jT3gG81N8Mveg
kg5KvzLGHR9ZhxVBvTwJUOXHcCdM9LACBONMWHnYQIq6oyW3ABI63qthU20OWxtX
BDqz2ar4Cph3SV4OtUqW8XwgG+emeaJpAVyx+/CXeM7hWORZ1m0Q6R8vBhz3pxIu
M/7srR6XsW9P2NAkGZxYHubaFygxmpuqyJqVz36CTlF+UtYrQbF1fkiZlSciZz4/
UqHqz1gcwpNz91DaTMXgENKcyKnOCenPWZa3mFS9tUPIqonSht1IKtdT+fvRgjPq
4uaDQuqliID2AVRaTptAo6spd56y/mup7vUxu1F/w/AGyVluA7I6BudynLj9TO/i
C36PHzoiEnaUuOtHEIbX7rQOWzaOj9Sko6ACYs8kkaAhwrP6UDSHciOwncvr/D84
YcGcyupovxabnkHlVs6O2sMfnk8t1MtZ4GVHPX7YNvqmSwRiCQWwBUQLfPFGjoSn
MD2zLpB52FRuMA+HmZ/oRRuvvI0llbUSZl1mxguCBY39Sx+4igEuxoN+0rHdahug
gKaLtcoRsa00WqkSFhD1kVX4/n8sxcVuLGa4f9DV54y0D5MZB/zqxU6xQd3uWvky
pStPv53yR5K99G0ln1+S6iZYcVxCxNbFM8SSPJSJmXQm814GVXhmQWFnU+2CaGSf
RBfwHI3hijyDIrgZBQ3MZGZA9FnjGoVz4K2b8uwfOrK11HTuwFEw43hhf15bmBe1
fxcPtREb/hiA0eu0gRxSH1z43A24oPhxFJKc0tFGI0B2mBwuSwh+8pajMqyAgbuY
0Ss30E0tkms2/ZjGJNB4qW1RufyTv1EKOSMe1eNT7747Zj0ymY4at2VgpgseQjMj
v+ha3rSg228JDuf6My4DRcHGi4JhsaIfIRLl5t6HVGpb95qWJ4whvgbLsRQyuEKx
aOavLcJECka556I0zVHg8OrwctWwXkZL4RIT1wIM8hDgM6zaQkK+1d55BlViJYLx
EcYM2aoseYSZ1nkSVDxmMe7lnEJ49ugBngBCjjSE68IVeBH1A3gECWge7uFU4nkq
+XoeuGKHE4tsHiG+mlPP7MeuHOZR0dzMJBJNUs3KBHB/ii1epAhJgAWvxuMXNEyX
Vihse5doHGwomGWN7llFCYSEWNLz3TwXs3WY5OJWjsG+gt9q5kYsYbLKRu3o/lx3
puLRwogvhf1o1D/YmaTdd5tNfUidXuLox/aTqhvOXkxXi6rl2e2Mf7yMoZ0RPH/T
FbFA8EPdyEu67QDOMC7mlrlEXR/il7uwVBy92fwEQQfTrVlVOF+YirxgiVRA3Vnc
BCjUOWtVn26jD5djUxKOHOTbnlqwn/99JjTxFbxqlYLn2DwWTSODlUh/sLWQnunX
eKvr2j6zebjjsfG2urSN4cfounl5KumZY5jRQ3rOeYqEszAx7f4vb8BwxZUjuvgK
6MmmfnH1hiFgSKCv33Qre6i1KV+vVZG2ICcoLv369H3mRW3Cc1tjpCWad7o8PmRC
sNPpkJ+DwYN/wk2do7uBcoyK9R/QF6DhP9xWuPwHrkbXLENI8uSpy+ObOBV0ay0E
RBlv8y+zNpRpEKFkIumkyPv2zXEL2FKxGpq333oEM0bOS5jNP9//92KuHkNn8NYW
GK59VGG1n1nkTdL4NEkxgoo0vIZz6dIuAe99aeF2T5SgQUvRfzSSlkYqVAaw0wIS
SfZ6hvoSmwTR5MuJ8sZlIman6YLysXE5ZLi3yJUWYi/DbYv/EpzdPrF/tQQwlt98
kXh3NgZIRT5xT01ER7uk1eLT6QFEA8gdOSES1+1Tf86nVvjiFgexPbZYxFSe7aq5
32/dkDvsXLjpJ5Ts0U8fgwRNWauwzLCfQSnT9Xv/Qrg2tlB50PdnTIhk0eW6Ek8b
hueNm+5EsC1Hzh16AumkezC/SpUG9tJr1X8aZdXHFjQDausHdG7MEOWNUMo9AyXs
DcHGsTaUJUXc4Py/3VvjfL3uolF7zLs8OfUlq71nygCc8vvCn2GE2Dkl9ukx4+YT
sc3SSu4jxCfvAbx1O580uP88aE8zr9sfq4wTRQmJZzqz4mdtS/JrIF8H0X8iqbAg
tjOV/v8NyNKfKEs7Cz0AI159DLN3Trpe5DHcFQVdKornrMHk1m2YzGO+ZxsS1jCy
czGuuIifJ+k+kBCHtONyUr7LFMnYyO70zzon9Qa1RVE2vAT2Oq9X9GINdWmyETAQ
yPcwxaMdlHNz0KS6HMTW2Xms+VuftBtxw4k9ZXtAzKR8FDUC6MAwtWHu8BYXzYtJ
nvh1tX5N/kIHy1CYj2OFJhatzDFkq9S+cBqL6uBd8GIUU4mIPL4tGEX/8WeGMt7t
ncBmFn5gntvefjF31zRrMUhCmfHtyH5XSYpCREP0clkTYr18FVDbQIKogGh6pOQv
aIIAofhAPsRjqVtcKYh29fQ+bzOksGQH+IMONL8GKBty5kPHAXDw5gJGY6CyMav6
nNRseqcVfsU+MeoHBzDCWJ8nq9V71P0ztCrw4vjxjLRttfF2+lDET4dHqfR+BpJm
ckrfdI+XaOON+agaLW51FiuSJBQAuh301/65u45Sv4kGCLqhOVZrb+y3GlXNFU2K
r9SS2RoIJ5XwXOeloCbEY9tFGNhH7L4NSSRqpaxLe/7MKzmSWFLSiLSSuRjusJ2C
AlT4rHBcSD3PQ0DSkLI5Zf2mS7EPUbXqf+VUiyR2pa8+UOdM/U9g/pMBVVQNhcBO
Q0d1O8nEb/Zua2Mb5NepL6EZ+GA8ue9DKJChkmK/iZEW4nASZN3wuKqlenIdiIRe
cHvxbhlNk+4ni+PaDYaNTNJwipj0rlsmHSIm26oCqnCEWumkUKAEQXxS3sS/WEUD
lVof7UjPf/Sn4nPPPEMcz5Ki+Pl2fRZ/dP73M8+O3YGMMsu5R49SVyvMihH2L4tS
7w7det+k89OoPlJNsvWKOuDuLGCNt74reAsnnIFET1CCWILaL941IekahiBFjeG9
tNSMjVhHOFSDA0RxRiPOXfix2ZxM+M/ROeSbThnXdTM9dYb1NokxYYWmdOv6OrzT
ZbblfuVuGofQ2M2+0yco8oKHfKEkJf3Gu2x0f1PqOpV7JQzlncZtE+thWNpXhYFi
bdCIOJuQFAiOCh/NZeUEad44QSC9YvnRWpZGi3gVGuRDQkM1AA/oF5cF12m5y1G0
UDY6vUwBqgNu3LSwuAZ28DNmXPkg1Ly3mYrzJiZbAgnME1ArlgkEJUG3iRvg93W1
bz6oXNuTno5Cfj0W01Kpm9O8zfx7AJNg/3KqC0CJPxjH/eQrmF5eLVq/RP5W2evt
GOxlaKYcRW0lVjG6ZHfHhD70/L86RMtL7ld0wHS5SI13uY9EqDTzHF8yD1a2gxuT
rs3NJMKyLFWqtWHKtFrbtCFihtIQKhd3mc+Mf+NGzDocudlhqTYB7Y0FHMoyQWfk
i7MCmSjWNvFluE9CrLvz2lvAAJSnFIV8xK8rnygxJSaZ9TnYP+YGb4+83Q07Xwcu
OQAGYVpS1knXFhD9SxIvJiKUkauOKbGNp8zey+svlGGUr6IRptRrWnd9/85mnapZ
AxtDzyc/nOc91xoaD8P17pBFOx4GPhjBGaA34klE0CLaB4nQnu04UHcDYHuT++Z6
uA01K6c5TQB8pcIx5NZkZGEISOOJ3NAzf8RT36Rq563PLkP+7gflDobpEKfIvhmh
SXEjHUIRorlJj724h3YSo6Yxx6pWWnRgIPnxeJ+QiXqiN8yTz09s1QMlsT2hv0iM
ECXZu5YP4SErlUB1GWgSEvVwqr8h285Ues2PByAie/VBxJjxZutF2h0mPKwErqQp
aUV+EhxHiwBrY6wd/91xhjMbE7sEYSGREiUHzqFnLBhGzAsy+KLqsLzlAmeakIaf
BLu6ndACmHE9a0ouSUrOGjj+IwT9nqDmB6A9wI+1X2zHSr0hB0XfGMwMpvCNS4sI
27jv8XF8zLqK86cL7kqfWtBM+4HGHyNIfL2KKsbVuKEjYOkCUHWm4TIHOKTcV9Nw
vByD95PmWowxJMIXryw5z2JL4OaouN+DIs1BqtdKscMSNKg51llnejK6NxGPy5Ay
u7s5Ev7yUkZd8csr2CJQSvN95+TJWouWIyRP38r2DTMz2fsgKJ/zhWPwWQnKhber
ubMaNRcgcYkLqV0V2CDslzGL/hC/sYdLYx2s9fODHM0NskgbTLsbs7M/xKR4FVJe
LARfsEy8Jy6mYc0hPBMKnmB+h5FtFhwk2hgsnPwJapajs2tpjDqK8JYHq2PgaQAa
CPQq54RSD6fdurSAnG+Jbe1KPIVtQRSnZN7VK0dThd8RE9LeE3vVHVyNNWetXljP
B2JKGow7URn/kO/qOvMDHFAgVLiQaB9i00JLTagPhnYyI7N51SkTH+0TwrSDODGF
wEC1TQFHq1kUwKxJHbHjfhGDSLgEjA3/BhpT4ZqHcvIWoQbG9pOYPXPqO8JtyFnh
sTViKHiOzstiIzm80yUI8jEdJ+njYZt8HBcXkDWgxnGAuyoMeDG6nOaDUEOpN3l6
pvsUG5dCLy5NVADkKHzKBcCp7t2r3u+008L6gZepMN2ySGsvVpde3GKBtDxoAITH
E58n6onF5B9v9X7o8IhED13tyMLnLJwXWPgsEPBmqftDsZt+DfQQ+2aJqV5Wj7ZU
Z8cLkngdaLdF1EXvwSBaMQ8bQ7P5KIRMn+vw70yn82Y1bD9X3SMyJhGWC50syk9C
hSFazIcdz8TzaI9DK5m3nxxRjKEqoMgk5sF8ANVzjTWq2uV81WFvlHDnQcZ6cN9X
ppn7bH97O9m8W5UbmiOnn6+NIvfBncQl6XiCip6tIbbXKdn0NJfZ4WEdeRbSQ9HT
/Gvs0oslepXuoQEKueIdCFFrA3cbL1ZuJmElVXL0VNfCbgkfnE2KRMLudJG17McW
mE4X1zfmmHlROQHyQbMmD1E0rBeeace1NoTqMZXJOXXiucAaiy2uf1LPNMyzgyHW
dt5OgHuFWz/Wrh7vKrYAKTH4GDQxz4U74m1H2uYpXBSCZmnqZ0Ap7DpTAZ9O/KCK
Q5KNn4glxl6ZTXmDPv2qN4wbVq+xVWoZ6jUs8glZWXfI4ooDHqrKjVjNr8+a9WFk
fGS/1xprfq1HoNXEP45Pm0/RuIxswWOqv7AyXX/5JlfJ0zG+hVS/n4VMaEJMKAji
c2SfjzBxq5Ur54BnKN4o8mj6UuR19v5PTofYKXAbXlTClUnJ5Oq67TG4Bty3BUfl
mUUk4WlUEmZufwdUZYWLwUJ3b/FdyqBEILAdcf8unPpuxuN2BX6JUBtVn1MTGq2/
vJO93khBFB9lCnbfmoN5QHrdfwvCc1IxWefFn9SXSNn8UUanuspPoeMNlIhpjxf8
W7sj0raAhD3Y1+3x6oDRzWrf84PvHMbrO875AwZAQjzQLYca66k+DaGXmYlDREPp
F29e9L1pD5tsbtLy71cVtKgye9fUkQKNahPIJjKYOk/ZwK4Pmzm7gUPWt4C5byOV
xeiV0/GQUcmYvXn2Uy8nnGDiEojd1G/gYgp1Ys86SpVzr9OQVZvB3MYEpIbUs3ji
9IN4mYxK9UgrEN5zoNPN82YQczP7XSzBdEUC4Ph/eUApvMJOi2Y/ttQ+XAsU7lwC
ViNMfVme+dmzQuFZ0dRQEqZF8/vSHwaANJm1471MZTj4hgbj5EGGkHc6D4stbF7W
67NnHgqaAgnAxxykXNHtWtSF1CyD7X4GRAN60Gdr1Q2Avgbb/yLvhldzmS2KJI1V
t6aRpjezo2NAIm/y7pen5hAfSljmBwHmZeJiS6qpQFivLzfslS/K8fqjh3d3cQZZ
5K80f/nt8MQE6fbfblP9S2j+OOCiFSGK7M9tMF9Re2LkMy5/sM5jkrIqC8+/Ya6V
9vu/LMxnM67/744D34nXeIj4BqsUaTGHQwNFL+W8eqb5dJBedu+V6SYCLlxctfRU
7/T5oNIhlm63vES+Px4eJsX4Wyb+6YOzJoYyHWRHxTsnDKrju2+8Ddn2b6BWzQjD
tBO+zP0k7oOTH1A8uYXqjdBJ5QNwOi9FQilUWktoaIsy1RK68g3BgQgO9JGXGf8H
0UwEjjafhINUF8L3SxHO3mnB2aPRfqMXiQ88S16OS8z7hc8f/kNFcEr25yLlWFIm
62Ot9JRGjmVDrnCtqtEaElAD0kyPvPxKlKlLKjjUFxboqjafHFNACCScuOsmB/Lr
rTlxil8LWdt6RX8TgYDZh2pp5Kd4ZYYvUqNwJ6Ho4XfeeTPZhnwsgD66iMvKa9JJ
CEBw9NMe8r36RtbSDvU/1K7lfOnxBdKkRbaTSnt9Knf6ssNUCiEyrq+ubO1BoIAV
q+6IVCzqqSWdzV4d/cKBb2tN/dgCuxyVxX5N+IM4QS3O5anyyxEhRiL9BYTsdBAF
g8jHMHv4HIN/9kqWdpWqBgBA/KiV0TIs4D4rl0JxfkP/A8ydXF17jzHiVi9NCVsL
35h4nj6UJT+8vK9isvZdyw3ahTHqWkZsHPbukjQfsWwVrOvWZMvEOqlYSGiVWo8J
NjA7MwNUQUSJrT8PlcpXeje5oB5krNTifBSeEyctHJHARD95HmzjUoWWDJs2x6Q3
BTLX46VdyMBv5SeW+1NHQSd8UrRjVuIlqgVxth8e6ZCj96QGHe/FjhV/VIp5+xxA
xn2lPcnS0lrWjgF/8IEyEfZhFhs/F4bQkMCnVaLOJThQK0fchiLP+sh89pk7c8nc
XgIRc/tg7L4U0/7eRO2v48VWsdl5VW/pOvzb3R380COvn3SBDwUqZtyVbV8Rikq1
TfTDJfIovcqeQOihIbAmMW0/bexfao74qDSyRjdR5qskZG6O6YYmO74aXdAaiYkX
dxE6W+eulQoiPJa+idCtV02Bhmc7EXg3wQRg+YEwjVzyaFLPSFcbo/VrFu1hi1J5
dbCcvPrSCTyV+xigxK3M6WDogDtAns/sxe4sNSbamWPVT+Zfqrc2gtX3k8K8sbLg
zCAVdLx0N7TjPTreBfCErFviUTNl4wYcmrY7YuvYIJYllAUGuWGvjLrrO7VkC6jQ
WUCcpcy64gUBWiCG4QVEf6hDRdj8Vw+3wlY09QYMe8AqyXvK6f1sAncz4GohxIzY
mfAA9MvC5kP8cfeykfWmFU1GJpvqtUiKdHq7mMJBdnDeckRw77pMWwwmkrFVJoVZ
Foy4opgFgGlTHGAs3Vb29rdkpIf5gYzyK4fK5hU3IO0PiW65A8RgCd+nz6HtgXon
bz/hSCjYRSuj1da7EWfY7tm/FQB/XhTAfRoxRVDChapi5LARX1DDRwYpVDR8WRME
37y/TgQOkHnzdSZ3snYaNEHfGy81/89BecmnpY0z2c2ocSJbvv3bjkuPm6kkAaEs
87yEd4HMNA7JmeA80uYPaUc8/N0WwrxPLKTvE+6VmLT9BSnjIQbmN3zBXISTnguK
i9s3K3tlQy/C6/8XOAQLZKXclnZhJ4kh3BTl7A2pjyXkZFUXY/nxCORuEJi3wJEU
p5o6jTcJwbiwlgfmSnQuA9+M8Jpvog32iZHG3rvJfc+S5nJtiNEdOs62FUHqdw3l
svanGSLj+aUdVoF+Sofhd7CXRJO+niJ/s4sBHi0lMUvYqJiG9r6a6mS57HwdT4v4
obD40ihqZkek4EPrupuiTjdJighu4B90JtSNaO7rDrqLO8OpEDc6Lu9xZvesc0Qk
ioy5D6B6CK6uDS46y4/ZyvY1sASJegGhgUEATYYe93gwyvKNWMlw5clOaj8VvXDq
oq4HhN0GwWt/PE7NGUNBfuI9RpzG3xn4jYXXhcSz2ZQUEI+rMQbjSkELLIVp76he
EGC17ru4zf9GBLJlfAM3grp2QZfEQMw4xtn8g7qtxOOfHS1mKqcV2YS9mQeg1eZ2
RLPgNPvN6Yzx7vmqIwc0Bk8ks8GAJqyYmpIZCs4xXgDaM5/lzuwmQGS13UbgOsH+
7Dg8J+vd7y5i5zjDito9Dfzg7GipMQJvhGES0xXWVs2PQ/eakmdbf8G2XeAWuNsw
6IUy+FPchmAwAl7WOrgAIO63gwl6KJhS4Nih9KPP1Gm3oItTzgw9s/BSdxICwHLW
9dY4ec8L696022GiWToMXYD+s8ZgPildx6aA1NrDxX9Fuu868wPgzF4ZtMJtTUXY
2kGTRlNoUdFM8LG3vu0bwNh/3x/fmgGqCcRzQFWffWQ8RmHzD1lKXl/fFYUKOmdB
o4WqnLG4WUKuJRW4gjF9CcPXZon/Vh7F3B0p+RUvvhdj1g2BFZBjo9NpK/ivZ8yB
TKPDb6O7AjT2DEM1YLgzNKof+FMIpbnHeOmtt64CVTzGEeec4XoamoT2f3HBf7M7
ywRwEVOX4YUk2R+I61VCdrHZF6kbFf29Tom3pD8o5x9NjwTwCMvTxJbWXoyKeBrz
5jlwpogPcCtjWJ+sIvowrIJn44uNATPHMS//ZM1lKXhERc2Gew66Gn7eU/GYKOI/
y4G+thQ2lqVXTLjJFJ+OaG7LIEsfhV/yAvG+bglmeQu5r5ifnoi2V6F2G3vsmPuQ
oRRUDTuPlO+ElzpmU/E88FsPDAL9zL+3lu7zRNG/RcLJQIB1gup3iTm3M2iQxUfU
KN5kchE3OHXy/O2vAUyHeC3Q/Xfd0G0A0faoKT8EwtRQo1fujxqUC/tmgPGOyrgU
rb34DdnQYT+H0rMR5PKHeSLtX7hcUjwKeIcx3G622Be7GV9/KSFBFpnDAqVzdwvw
o8oBcxBkblHXvrOCr6KR41XUhU8YCAj2q1PHtHrD+Sanh5GPXIEwsNzzltjSymz+
MppseC2WdiF4uWQTczxifaT+REY/A9QEUdiQsIBhNrnUFnroLoEdxeyXwXmau0Cy
Yg8P6W43PHWKVUUSC5xyhfr4ggKN9MMQGzI7MgLuZtHXiO87Bi7yVYnl75DYzH+E
1gw42Eo4slZKIDjGS+zW7sDEom5XkDwXp1uTZyBSrCbXc+FdYYvUefbUMbo8Ykkh
r/HMf3ivwK65fYkgkW825kKufFmwx1YRhy+eJi/lhUd/m4e8gvcbz9KTULGHlLHh
0aVUyl469kQBeLN0yZ5Sw36/oanEjELiWtIR+hQ2ygG+/aJZh2r2BcKio6v/Ivlx
dEk8Xg7CbT03+R/ee8cCdv4bL/S7hlgwpyYVSsBmlsoJMIrCczVHt3E/fLTTztP7
mGfbbvOzIVXiBqd4vkci3LIPwsmr3j4u+jG0hO6vf+BXaAagVJKZlfAmdbw175jR
np0rqquwwzFDGwkARmTddJ3WNQU+1NhXSe8z8oI84xdE4ohd+P7lUpVVAv5TbXLT
6iKKSkFaTZ1FE7sYdtpZebAQ3BhKDMlx5EFjIM7fxGWm/6sYROpSdZN3lNoFtZoU
TanXCmAYiQcRrnKMujvg0qhvdp97WM8BNfXIWOuNxJ1HQirFEJ57Bd6OSfOdiuMs
3FWIxqCW/cGzSuENaByaDzozROx6vb/zxqk8vThyDGhkcD4vrbdImms5hMWz0R8H
mH/4l79IUqP1vzI4Optc+Q6MF4bHr1amLdU+Uvyzo1x457UOyWDy7CYV7toZN802
nP3LhwRo4S2k0wR3c/AE2rbuoSckYJMIltncmJpcpS1Y/U2AG1ZrcorWPjpAZoix
yNz0c0v42DryqaxBR8HtShTAAaHik5FQuyS+2ThWgk8TC5NCPfMNdUfB0BpIm5Cg
AI1CT9m9p+/ryU0zuW9s9uYMNaaMa7q3KDdrSGmMNL2aJxQxm47MG9gjICvnROXm
vgMWPC+zexwXwrghDmxWOG7ZLChlCwYWth4Tgqx2I2Yfsr71QjqVn7nxH5X3MK+l
VLkx7ny8cB2e74+86PtiACuVwNMP2B/Z/HmxiMMGqwf7Py0PKBMuzhdH7AlmithS
tbq5c5+5NE8nbmszaLgMTb6mILVha4hYgMffIWO5vNmSUVhPFmjVafopQYSxyzva
3VseeFYbUiQPfHK41hIaevtoIUey0nmThXz413lq9uZRyzk/3orEWjKZCrdMBxPS
9DN2l/VxL2T/A+IMhOjYgMtL3whXRRVrFLzoBAFEjsxevaUvdBXKbmz7zaodQkEq
HNBuksiYgRBREIQIHjYd09URdCsCm4PcbI1UCt0MvUYlkLqm81f9EHApbwMNnkgi
yh0xceM/nyji7VAlzZq5ZWthcWGSCjq93ZeyQH0ywA06CmdIf3V41TF3enmAFEAS
WgP2tvJP/2DbQfWmyg+V8MypjLTsGmCmiuDbvStAPS3ANPECDj7zz2gBAo0bCIFe
kpkxui6c4av/vzBgzfcZgY25M34mqajkC9wqfTHU5k27tn1D5KyhsiT/sULQMKa2
azZ6owtyeNdVd9OHfFt5F/4tdzgsgbhQMvUw6rICmwML0GQTp0xj3eogu2DVc2iN
ccagrqjPMQBSPlzV6Na7lhTCDZf6WIoB9+dvpSth92jcNHR0VyDZxb1NfmHmsV22
MJb/4TqSRmsKqXyiERP+EeVs4Xik9n5UKLBRjzdKyu3NI3HBIadsB9ZiCXyqNSrt
57mBKUV24uJ2li7x9aSA/pdrAafNSDtw4u5Aey4i6KwOVBwvar8X5nwqV/i313bs
YCo6f52PkD/rkvd/4xG0L4Z0F+3LeQHIKocsnrJH7/ABksicv6MqeW3pBaP6VGkd
v8k9OaWw1wrO3SfX/F2URtCCVW4WhJLDBN+o4PiV+tIjKOaaOAp64RAaioxJZ+QH
JHjAUHb+qbIml55v+wRfxTVwJ+jqfUhballKgF+ViW0gyR9upWcjOv6d5E28+BnO
jKOtH7mInOkYkUYymOA03iGnxBjXq7aXWUJQ4y05ojWna4ffG9TUtwyXG5vnBlry
mKjwZ9RD/M+V7Zvhxb70H754eUqDLMXObl6G/IrPstVV088bFv4Cmk71zPl6dm3N
Orq28LWbGQB/u329QvOy6nuCtNamg70TLCJtuyjq6CqE4D4Z7e2LYgNEX9Lugiud
+EsNeAOneWshFw0XBvcnE334CV9qkk9Xs14UWfDyDor9R3U2Horldut6qdymyv3q
/9+cyz7/sbrlBQQ4JQ8IuLCw9R/j+RM1w/XeiBna33Y1pNVD9uixk47YFREM3jDv
C02g31ifv17vveLYbLf5+Q8mXNmsd5/uzHgky7PFtFkDjwCIOqeEkot2mIh2jxLI
6amgvhkYudaJ7X7vBPIKLKPmXJyNs49rjn8QQpE69Uw07fNOPLdopsKrxJT2WhvC
DigLyy7ZNuK0QjD8Jomqj85d/lL4+SWsz8JbgpYHHiFvSCUmdbYZxOuhS+6Y2WKR
9Cx4zycawAXmR5HB82k8CyoQkkSVDYQNqQTVetbcZO1tEHm2V6CSM9usnbj0zed8
oqKaRCDQM4pD8Nl3eV+NMOyiRILMjA63jbr3To6lQeqIusFOQLZxV3THqLjd4+ye
mTpzKre1UI1uKZ60wOEobhiWEkS2ytacKu4fMVLurtKA6bTSk9Zxl7D5TSHt5M3/
e6vk5CdDqn0U+9q7PVatczrK9qgQ2VMnCN4lWrXRLUv4P/bjZjgSxMetX7QRIq+I
2dvcrmA2SFDPd/zfdI3xEuMFLCSEVCfacUVwLR5bqIlh9sU7kj/s+FNAoeszWzuj
TI3NHn2pgqP3XXcOWX7Tean7NcRuQrLNlaZne4T/8YsyRBMi/tGHlfhVw9oyo75q
bA4XQSu7xN9aDUpNa4CP6x/118z3mRnxZdiO08DiDWk63+WGr52JH1QrZWRbKOlj
nzJEl/vTCsyH0K8a3LP6tGq437ZCB4guUBSKfYpqezmNQwC8pJgYClZeGPJN0PuY
hleSeMl6wa9xBNICeE1+s7Ft030jQzuuzgsN1O7TbtggGfpa2ntFQsi1PD6qDnpR
gJuhZfki17a8rddOv+fjkJB9Qp1FRw0vyzfT8N23GzeSDgkNhpxRKI6VP9J3i+ib
gg8rPj8Ipen/5NcSFCqsWBRVRkzgtcRCu6KWzJLKXZcmCuBmXNHw1G/lGvNmGw56
ZgvnNkQRHpodrzsZaotm52svt9y3oDt5HXhBn8+0FyF0FFH0JPmrkNRCA9i1GDdv
iyjqDW5FObWEgxy2edrg4YcASzfCZMbFV+jLmaNcD9DFLsrtlQ+d6DsDBsBq1FQO
gGKqHU+9amxlEpe/ytfyFCh+Lr+GnFe5T33JvTxBvksKWUTizkuJdb43jSrk9mxV
E7TqU5IhVEEIfKE5isBwctE+uP5zY1cwagRXlvJ8ITfz1/4fqgM5oy5kkuiUPvLm
yJxCuH/5toeJ5lmCh1pmDxf+YS7R4rLbEt5yeUrdwQofju1sUVBba8Zi89Yn0gcR
jnbhw+8TNFJoTIFCB3Wf4kf5Vc64P6ysIAj0MFB8sxkV2l1pR1L4Scy31Cmd8fkd
87Vbp5beJS68k6gdoMzwQzWUcqTgGMB/MlD6bI2Zkb01+m2N7k7JaA1dn07S/Rg0
CZj2IkLQEy0LiGaSUgnrH7GdY4vqRORwVW7bgRL/MDLpny+Y9N0mTdwUHw4smqHP
NW3HXg8PTW0jdzoqUCGeliHzfyQUc5fGyrDtsiAfnIKwCVPBZdSPG7tsHFqNuXfn
UgbxPylgjZQOLVsqiMgZFk5ze41XTPUXsl+xmw6D5sVHtGQoduREQx5PJcp1W+Xj
pz2e0FDK9JkziFMxcyxfx/wncE0v68NEczNljs1XlY/mMc1gc6ESBOKk3ZiOy2Qv
gu+xNY1kKf38FaffzotUul/2HzROiRYa8KRGGF6PXitIUPM3fCFbeSKcfX6NZfrs
IBiRK8ubBc3Xfmii4ytmg9go9NWw5BsNozvk7Y08m2kS1JiYnAuMEQDU7RHwuKBx
NFZbB+Q0rpyyEwARXaXsuh8WagdaZiuz8zyHvd51Yhi2jqrvcyTrd+zASUH80GgG
oodIOpN3dh3z8Cv8a14SZNoOvx6CIegcYLpXhvLTHoqmnIf6tVre739pKUQbvDK3
oUYu24rkku7l45QQrA7ZTbe+Ebq7nE3O32zhe/A2fEtPGgAYZS+OCm+dW+ggeLzB
Pm1FS6iJElTucmK4RmOBCg3FL5Z/xhALJ1ry9exhYvt4QrDZOppurPoxj4mRJegY
WmIE1SJki1GBYs2hTaGEPkxxgHFqxWJUJq24GcMwCk2uenOeql5xthcGZ6rSeZ4t
RCpbpBV5wNnUmFi51+Ag7MTSXCLoHH54x3E6SDOKRRAJQ3Fmjc2G3yEtCzHh5ZD4
mjsYSMNc0m6hOU2NE2t4j9SZVx7GkhCRMr+p9HMB5E991aU7EOx6b28PPY8sMJc4
wT8awH1JCN7y6woFDIrmCUXmMyU3Gh/0+gDbOBPWAvoxpdu3CeW7o8jDuX9NKsGh
1CpE0myLosJamczt1x695grQeWiS2wIT3Xjb3vs0KeeKMnzylGh7QgS7yshKU4pt
AEfQTZphVtn6sO8v+cnU8TwtYT9dxveVgKieYGeeQTVH3lRe+McbRqkQKT3QKdFT
35Yg2DJQ3kIZJOo1XN903+6KDC42Xk0ORYW4Ia8ln/yi6hnuoWE5wnU0+TJqo0hX
VghnIO+aZmaSq8J243y0JDmHKGyAmsOTMULO0Dyx2yQNFXVQ2b0WTljO6iJ0pkya
eHh+xLDEJsXQu21x0wRjTaj5t2BgU4XghG+cHXhm3fPuzHweLw9KFn1IwE4hwntm
AqRnF0OvKp+vpPg7sId2BohegZpMRYz9RRbea1H3NHkH0MU9pMkrwMxcPKyS3897
RLnIwzFyUFa9/BUpoukDwKR9kxFQtNWSm/77GkIeFjK1NdQUlb6q63QgfnoWBk4k
e2BP5ETN373nqiqGVmPhkDKtChRHEhtMcZU6QBInJeGi8T+7vxF815S+2g7eHgbU
d6PLS04DvvpA8mlVF40zW6O/FUZg7IfHCVt1Lwlu0Bulsd2dCYTY9PKIR+R32CMf
CVrmCWsMCXFuYrtia4K8wBlIphAvz2oELsO5h9c0QWEMFvUfmfahcNdgCU+eC9c0
ESEhmf79/ZMPU3XNQydcXLYIVR2qeZqVGGlihd2CuB9iNUgxiqvRCiVomIJRijWR
j49rQQt4lhb81hKh1t17IyTbgmZMnYQzp/icLbYdCZmw/LS0YBms8ZJfScsstvbr
xyjm5zuD6XR/zxR/7tBnfCpyD7gUAa3/7qlMr3uZppCgvRBVfnxFsmeJ7Ygb4AVf
GBc6gw83T9Ro+RftypjldJ0JWx3LWW1ggG0++IYzdX29OATvmDX4XoQ7vLcJbIo9
Ww/WPtjXrK131KeogpHzy7aa8I5SunseD65CIy+CmOz/sLbTJ/TMu7ers7BNH8i4
wxLpgFKmm9wPEIWGdy0Xgly7zR+G7FaA9H3JA+tVmyoVNBv+9Jvg1619f7RAyQ6e
Ch6CiGdZh7KI4Gk/VKmAVuYndZbSfYjRtz04MIguxguUwaREbu7MJSpIzKPYq9zq
XGijIiWYIOql7uMs8FCbQAO2J48oMtGmQJitJbW/wiVs5uzzh3bYPxTyThQ3FtEE
WXlSpTHWHViw07dM7LlUAwQq9yWDPx7CuZ80iHJBIqzfZTLY52WMoX0W/qBsvymm
/Jsz15o4LnFaZ7ONWnTYjJuJv9ganCulj9Y3BR313z2JVD6HmgbpjPGFCf1tyXnx
mjiZot2ve2vUNTAbS/obu1sjn1PEYE6dve1xmasC4dRbcA/7TSDpc/qjZ5tgVajq
RYYVkHs7AxWGI5czygl7Tsm+JRevbXbKBYq2I0Lilwr4LQljS7ixjZw4CLqPf0mL
E0Yef6EdriQoXU1pYGFqXpJrDZZ2ubKBEML3F2lcayF+atfzOz3t2wkhG0ZpWm2N
qfxWRy31vKXv41qrhUewIFlbO+suhRH1KSBLFgn6jFcqVJegXG3ALpwaXWmtd/dr
plwdwmbMi/Ky3Dn46wozoOTHlxn2QqipWiSXEqEi2v7aD8x8+k0oeH7xvd2wSC+O
L6pLBhPYB72sWD+F0Ual69+LsqnQU8gB8Lg/AxZQ6134JPTu7fDnwWqezqH35N09
CeHSI6Q1azcX7Sqbg85gh3gKWx8739pV48LBI6n42ZfzlENnq/AuFnEZTv4SPrsi
HHsEt3kdrPlOqUdztG6h07iz2IyZKGaJi834N7SqIN+MB7X0/FlN65slsNZ7Z49X
1WDRP/xKnu/wqSAkcKODEUsA3qjW1r8e0aoUbf3OrBDS85cm893E15Lt0OwZJl2x
iFp/zKg09HUfchGAHbfACC4nbELagRRQjJl5rdJx2dwHscp6gcYv+GAIfM2ut6jk
s+VA1zqnzE/NnEl6tELYdSrlykhE+NMoNusBtKyu5YG16/qjPe4vLXSlaiFz/SxC
8ZqDqFGqfEF9E89eHla4j9IuOJ275/DUYvh78iGablJQw56XxHVDiQYok/KUKBlM
EozA6Ly69I7qz2ZdEKTn/fdyFsBwqlL80ObkxIVlX6bLT3sKloGLQQXJweneLj+m
yHIN7w7mXHmTq0a0rUFm98a6lrWwuBAKcLLAH8sImsZMW5nz589OoeOLw7KBRvmu
j9OgqSJKnarF4xkxPe6vk+iqOf9vZCy6AG7rQfnPyW9AgMKnmdTXwiS9kdJBIwv2
VRCSrtQcwP2xg0+8Olh+gCCgjlXN2nj6eUrCFXHA7VXrfmdR5mE3OKcVpnnbyp5D
Ocn+FPSCuhYJHmJL+K0Y8jCYMCiNUTqsWoIEaI3XPlJyr9nAgoRMpb8LxfMZaBe3
JoIgxCKNPu1GIA4FFjs54FcvMr34FkEWZ3gNV6I5mL1zDoBsd79ZitNcYlSkkO1J
rHsdT0xqlOowWfmwOfzNHmlxcD05U4vToUWl2Qr8gvjyS+jBR8XMNyeT6cBsqGQo
u0SsyFxe8KgNi3EaX84kPULgUf4bAxMs+h9Yvv1999NAXMDZ3kZ2DtYiTtsbyc46
gy2lGIwc2o+xuS41FjmQBX8tQ4r8ZjDW4OKjaM9uz/JRT1UeS95qmEbpZuUxcWI/
M9iw2z2KPCfCw7SXdwSVYsyaSCxzvrWfL9+rxhJKxy0cSySrAzdA3UYJNe0yjkXE
sBXR17rni3QILZdD2BSurSxCSfnS2ZtRT8sq/+0sv2a68SFC5kEEVKnEDi91KvZY
1xxu5wu5m3Mhwtoy/ppIC/K7O73n2DhBJBhICsHO88eil/L4CUAZWJBIybNfzroh
iObe/1oPeaW1LJsNVyWivn5Q6+Fg0tEXVYmvxEslOJOvB7TacfWm+aE1v18+Owcr
t+wyb74NBUUag9VJ9wWOWvtSI7qpoIT+KYGrQllAWR5irZS2TrKAbis+Muw9Af9w
TyT1AzOgJ0ALYvMn1suj9bGkD8jIjphQXLJ9OreWSQSiyIW5ibX0ydMZX7OU/Phm
bkmABKmNVDqTk59TJjVMXIPvI+r5vSv6enHiDxuVuV2I6vYeUln2I6Rs1VZ2VJB6
/cZncx/N/ZZFNkJtDi+/3dZ4ZFE7jyguQeZRMfHv8OlQqLBeieURe/rYpaF0YZpE
Ok7trsWkBg9mCd6Plzt3KMQ2oEfP/bkfDYcYI0mxJu2haG3heRZodn7iQlcPulO4
VI/M9E8U6iN8k9HZW7b9mRosIgch5D1Qy/CBYssbLVeCXg6cL6Bn7Tl4XsGAnWTs
wyOHI3aMlQURvf0NhIbDCzp5BcOk/HXEBw9+LEKe4VlCWbftBzKmfvz5r/yery8E
m/to1RqCeGxvJ1Gh4G+Pjc2CfQzxT9eVJq9+APZaRkwYpeKuPrO2Smg5zT3oE6qO
mHazin2T9PqCT2OOnQtXVhrlAFbCTA6dzr8Fda/5VsBn2YqQyISglTgIgvcB/QKS
LBHul8yeVeSITcBVO6FBLjl5L55zD0YxIxIVIPvauRDchzCoFpRoLH1mf02+B2wl
G6Oz1L06zLNi+n6c1FJFX72ZN4MWpt9bsKDHrGwrdRUHQT2DCcE4pSVfCnuGE3Bt
pFmeaizcgJgg7su9NsMLfMW23xPylHQ74OuEOr2LeF2ya7OyRA4yiLEzHp7nR2kn
xpu3zutfWn3Ba/1NUu0q9yg/2e3QiZjy9yLBHorlYIT1efi7SSUxBT5bRfKeGzTt
1PoHqOGuYK+puVZR/73dsK8h8eDXkoH+OrzWw1ixjmZ1wtBR5QE0OE1nC+Hdi0Xj
7uLQ3i/KL4Miq5JcPcWBmk9FppGnmXrOt0wT4NidPdaBUZrbFM1h28QZ2TNR2QLm
VWDU0uvzyBir7b7gBRoeF1Jmdy4ji4R7qIUHkaKiPaWuHliIvFOE+8z8h/r62vt+
8dirDA7h4vjnwgwYo8yqLKhq6Iye4b1rPezH0q5GsFrdp7d2JRIQJMtdPj8L4fq+
d5FS0q9Drs229rbd0KUBgl85ugZGt8h9x9VGNVZizCHhYvMMFxuU6W6wwNKVqewl
LNRwgKw6wJy4zPYHKoOOCADvyqAnXhcgYoMWO20tjrkGSgPdQprL7FihArXSPGua
RAqh88+i+g4L+zP77K5WoPT3O1gnXNtIrgv1eEfpapWpk1+MnYUs0ZKqKbJs06Di
3Q1o8JfMog7y+VmWBf6Z/Ze1zaHqpPi5rSlBLEoJrndXNP8RK/SnHeueYWat0Rhx
xGBcGyK4SobqzQ6YoA4zK77Aq5n7z1zdshwZFrRkpYMi4WrCZjhnGA8cV7UFqZqO
OvJqKn0XuWRw4nQMwe0K+OiIMhJcrbquXlXtk22MpCu09w3/MD5gcPz57RzP5cbE
jGNmWMi7i0neznTIT7bwhtIXe+MblsDUfYrmqUtIE5ChmL6zNdSyWSfP6mMazwBG
ABLHzGSLtFOgYagJGJSYNfCXUAa+OSJ44XN9Udvla+m+L34OFmmvv5C7BHBmVsm1
VDGAR0ccZtLfKOKDD4q0ujlQMO38DzBIiGMOQMCgBI/xuRtBBWvKO3kDHCYN1WXI
Aya2pW5YXnyHpz82oOGaolNLfzaK7yDfuKVlPCnaZffJyE89k7r2dSI2Ac6JfP1Z
p5ldDhnFWOUs+XFYIhfxpaPR0sANf2Juvu8OcswdFXfoMgyLoKze9N4wFouvxdD8
NC54w1YQbM8wEvm8c4A366zZOSa+V6d0zoFtgYWJSSxVKVk1qSVniiXYY3q3RE5X
UYDHNdN3nxF1RQZd+o3cLKFSKF165qFVFzXuZG+i0qm7sJjBEp5T2KG4joWr0rJB
ZxLgbqma13dTg6Vy9IhkA/19AvI90tF2KknOyhWXe7xtd9b4+2u+pd8N1hHnA73+
OgRlyR4PzywlMjnh1svzFq9+4czejgFfT8kQ31jiHBi16J4kTBZJVNHvdVciS0Xp
xNiiAxYghg6xbvDRMdG8h/yPXW7Csq89udSXltZfP8v2eG3TxPI9w/x17JSzWXW1
xxuoR7IPUt1ghLygRFFU9AOsBHdBZiH0rVQqZeVMzaq5Jn+r+jIP2rZ8Itsyrs2g
N//q7Zcyaf97xutCbBxly+WKuZGfOFmuAocoI/f41oB7f76rkQ4jilvJ9ifgo+OR
foUamHpHofZm5s8eeJkUOo183MdCy/vqnKr/ra1hJZPFUTOr7gGeqWfIuLpBzq90
bTD1G+eEaqJellHt+U0CUimv3kDSIBjtV/5hzjdDtbm8ZswJ+Pz0qAt2LP2qMYlM
0NjAXWsFfeVqV2JsPWhmMjT5p71Wr0fDY7JJoh2Gh9f2IdPVdJV4c3kB3leD2R0O
ZmZOQGz7ByHCX9P0FllPNGuPCqpWhlPnPGYpLZuruR2ZSIY8fAg8dxkPZA0PtxGp
1OnDRVVcVZq0Byd8YH3RzL8+ewmmIWkHKlDiAGHfqppfis57UNDSZNhmhiHBTbq3
Ybws/wAORQCpZk6nkmfXeUAQuCaZ+Wzvo3VPh/jkfC2D6vMBfQ7r4jFeR8PWwXMO
R4DoFVr4R6Zd//RK6lKWfhecIsx6MDhbZO6WEKxuH0liK1kMOYKxEoctWP5wJE5O
qwODXscEGdoXeGLu1rnHzDVDE5XJTNBU9HDayqGPI7JFEJL4TwuYj+Mb4qvnLK/C
2q1kv9iNUG/An6fYH5K9Xs5/wmzxKwoSimykE2dFKQmQNDc5bwORicdAqjxrqBzd
VTnWxSmwxCSaZHfvOVdkpWN8H3batkynUDQhTpRDi+oZXmZFk6WAsQhCQWhGtUXt
rNyTZ2u6+IMfy0n8TM0UYVGJZEzphqPyZnpC+ZxuUizlVAhvS99zKMD631N5riP+
eX0YllIadt/qbPudrebIl8wiBc3OQbc6sm+VUttgRm0oopA59BUpFhpPPH3Gipwf
hNST7MUISjgjbKF+UmZr7Jguv/AUfFo7x0xe2FGLZUMzfkcezJ00sz7mUHYdIJqg
9jiJJQ12W6umHiwcCtU0+iXU9RwbjJM5/Qh5I+JkOzf8oAfixIreFO6p/34UXV6A
VwNfe30Vm25NQ5QPbjv/EPcDn1L7qQ/OHbORgX4GYDSU6XGFDNUbPI4RghnyIhQq
bYFmLWRcKa7FKZdwFAHxsqTaMu2PuwEmTQ/zg1V6MqmbjrWOtNl0tdZ/DKNszFIc
Ratm2lFk1i9g1BrpbfAERt5KUHqerVgfbaZznsWuyrguDXoWOSeNQWu0w8Hgeh11
IBXLXDsEBjwE2Vucw5N+m266mqRD7ojylmVTr9DhlMvaF4xeki4JgexyNW3lfjrJ
Rfl2tBGMTF9M3WSZWBlpeobiwNe60xxm/iwpzPCAbuRn8em2efR0kAa8Om1N8cEE
BzRJNNYuXEJHdLM6HjVFnZv7HyXBzO6EluEcfYV5DjWXV70BrPz5/mG4tyLWR/ZY
c7g14WcYwFMjnb33yJJr+hxCsN/NqQ7w5u2RoQmccw8BCmyqFV2vb3TZf7OYnyJ+
OUr81p+Qx9vPrxK9BI8ncI88weVSi1HqM1EFk69T2Of05rEM/PVH8Im2OwJu5Gay
YSn8ru6JoiDPeph1GvlWSJ85zfduFuLbatIYzs3kNG7uzoxbgiLTJ2zqF1TQdlob
A3Ywz/2LQUGYCY0XBsBTQJS3WCRMPPk8tWsDrMv3lNzfKT0NxRFQMV9OGITlCH6a
08mp6YW2BveBOFpWH1Jv3pDgracfTwVipEkhRkG71+CD4nJRSxNFmPO0zCEfJ/O3
6/kTfKffWxb2ZaefB2LBA7e4HXzIf3RjYK9Cybr5ZPnVUE2s8+2dx6WmhKoEvW0g
SWnNjFD37AOQpXzvqcj9Jlgt93X8cbWv9E3ZbHsxpSi5DNbvtyi8r+1kk7Ci0Pgf
yw41RmkDZrnO3TbdIUND7xiA3pHABzEZWRvzsIj03/zlA460qTeHzj1PR+4KgFvy
5uUaUc5E/H4JfRNDmrdrPHiFKeR375wyBYj1GzrLvkxOxAcs868IDkalQauhV4BP
TDXkVk2VA5A/YyB/M6vojIEPxJPXVE14uM7leLzBDJpt7TWLxCCBefi/cZt9k4+w
RxmILL4QTrW+IIRjAS0oWYNeTYQ5d+VAyugFKrNo+tVSo9qOeCkNrXXmznuLpIwK
jPgtysRGiydJWJErccvSjr+VxOpj0Kj5qc/ZEgPV+fi/gUyesM9PJt3k3mkZZKnN
2pjoK49Ypf1Q1zap3Kd5EU5RpmnTy9wjWo/fpQj4HkD8hhBDo+R+qghMToJC8bg+
bCjtxTMayzbWKN5yLdfpJWpT9Y+1VufCBtpvW5afG2BisQqAbPXMqfJV+fGa5s3e
6B5PZalNwDMBwqlSFjQs8eZ6VlQ6U/rtPh/Q/FBMBJVaMJLqcwqbGaFgUgUyljey
jKY4syHkM7HKfE4dxx33iDbVdenFyW1fPR9HU5UuztDeuOxvXrlSVURCbNOEmQt5
C2kgWwaRXYg5Jsp+RlcPVptggJ7noNt4ryZVCgL43TcVP1A1FTm4+Yhm1qeP2w1Q
LV0Z4Tl0KYY+ejggCMVDSw8r99vqy3qPKVWAn0E0mwDOJCAJZhzgHskniaHIzYSq
Hrdrce2QCvP+dWpVJXFSyiSAFrMey7CezLzowDlUahjflocZYIsJeskJ7mdJ3jx7
lSy0WdWKYNjfyESrge28si3jRTskVr3cuYAosCvpIj0PExvC3yjFhcInY+qlD/Pt
6gWb+26HgvX5f1jrtZXhBZv1ErsrSn8I4NU/wP2nPpgI3UDLxZ0ERuBuGMYTIcYM
LBpcKsosEaEQLVa3hu5ARKKcx0xZrDS2ff0Lcw8Eof02GRRJkYd8gTKzT2PAvAa1
iUkC4wzjD27L2JJd4IIdB0fhyPKGlnNKSoNOMW9ph8JUPI0fDBA5gVhysPljwoWP
K9ycJ9MsjZIgAwirrB775LsCw36+C/EOMy7Eobw0by1an/4DzoUK4HQ8R2Bze0LV
FXxKyXctLn/aFmTYH0/pFCzLZc50S6MgnOJz7H/CWvM+HYmEZzZfCC4JS2uXsPq+
vVMy/C7vP6FQVxZfMKnTpyM/HsKbzr9y4XyJzn0gSCU3o9HIbmZHJxjBfmXd3tSN
JzI5yoO9ETapjucqwunQvOi2/PG1Ucifh/BbacBBafrR+tP8e6bUnpETYf8gqTJK
z+KMhZKqRmsmH+HUbHGKH2FG1kUlJKkMmjLtLZZ8uVmz9j2gO9JLj/7kOU63E/Rf
Vz4c0vRloenGJDSdtx9B/MMT7BvwhvldGhHUwvGo85d4ZN7yIfk4+A8fiE8Qj1oe
V4hwTRNyjq665TAf/ExXgJsymxkTIYxKGwp6XCUl5z4FLIPgn7ZGwJmAr9l1PBa4
cMi1jqrEDIkvxi7bSI3j9ey2XOBDSRwZmrS4jeE9rn8Ygvhm5GuWRAKEGZBicupW
6Ezo3XYOMnlBF0g/9hPgN+1+62t+L+kyTQpS/sfnZZJw6wCtpqJIyW3YY53jS3CZ
IjxaFZ3/9NhtCa1QZyRjawbadzR5ZSK8JGTNptPnOksWvfw5zNcUlJzYNWh+o59f
iUJmNaKl9PZLeSage2aZoWBeHWBxMw1E3vUZGw/vyXftfiBV20waP5fXTz7/9Tn+
AU7WN3ePSOTbsmb3SBZ/Xm6VkoY5ufMvMdTgKXUjQ1tNbCoLQlxhegAgiVDd/vC7
0dludBkg2v2iJg+Fa/FtJZ4BUDbTn4Y0+hCK3KpEWjHFdTTco8gZReS1soVMqBn9
FeoEu2DShEBTYbZfgFqlxCrbIldCS9ETNMIvvVANJDbUdxKeJ1JsP8bZlbTRQ/Xn
bONmAlN0WzcMyoQYTNNqMc2qddoIbDArcSwCt1FKwuxzm4uQzEe1hoOjLDRzjKgg
00HdFrshUzTN1A2qX871+0pM3J4qnLB5rxmsIlsfFCPuxZRtY219kZ+SjPljAbV2
j4MklFn10iSq24F0w21UavNOAi5TOVe0UpUXcvhhnlbUIU33MaQ+eoxOdB9C+6nQ
sfXVqqmt2gUAZbV65z+nPiPjNRykdFRjA+d81d4uQ6wsU26DLcV/v9Ik6UvB9U+7
98PtP1aJuckhBP1VBG83cGK1Lq0iQjQNR9T5f70gZQ9IOIglqTYToMALUhuk8kMD
pcYQq4P0olVhywJOomtKponHoOtFRexnE2OM+Gc597NyW8EKkUqicIilJf16hnqZ
Xy7yEhXldmL/B9lpgZjPmISt7vkYcOaL4/XBedwjDN55KrzN3q2DQxGGkwPFAhod
0LZJx1NZzxymHcHNw6y5OBbdsbHwTR0Xh+fg+Cic/WZPyd9TJFvvWQW6Z0CW20fj
I4UliCBUyqPfim9GLnjYKYYWZM/IrVyODv3LNpNJgwR5L9v5l1P+9I01AQweL6DF
69YlGwKLll+JidhupOflRHq/lWciUh6jL0z0fClrwqeWuTEBCvjKZA87Wnb/q5ca
sGXTjb6/qX/jHbJ8ibC/rcyN6ZRCSGj9df2lmAzF2Nql7xYEbmHQvEsQAywFjC3s
HpAme4vJWbWK9ZxNcjSodhss3I+cpWEu2qi3R/cN2hKui7TcSv5RgJZMoPt8xYeV
oe8+6jFbCO5AamSd8/VTLDYefKOX8dfuFC/yfEU/Tz3EUgeM2WRIs4+FB+F9G4/C
RL+Aw7eWm2callNbK2gsSW8Xd7xjTgjxFKXXZOFsndyeh8uZxFFp8hRLiUbg2Vdc
m7GvvVXiMKkxDHtwE4OoEBf2CHs1LPpOre99r0ElM8P26RR2V04APm69iNuSSPm0
w9ZjApDPveyYrAnKGngvrUhZeZP1BKRx+tZXPxJ+bKIrlNoDnv3Ms4iCnvozh+HQ
rKJwLhIKWKArwAkOLUhvHM5Kj+/ixMfWq1uFju96//rliszYBr+8xiV4fatP/p9n
CjgYytj7TSm9To83vLSrtRubvwmqcHzToYU6TvPv4wrNb6ToLMDFyWIf1CjUKFe8
/8Xc1Hjg6rvu0ZWXlVgApQnw2X6AbJdn6pRtTCsHu0kf9jlnZaaNuderrGr076ku
l7TjO7aKc6HYs/FAxBkq09SHL2rwcUV6/6NBkn3CGnfJULJ3UJEzGvBMt0GqvAJv
P+MT9A/DMpvqg2kOOVCp4GYM74Odez3aleEZCScErhDRjJRIHz9N8cBlbVmJvyl8
xG79oSu0TWyy5gGj0lVW6WIvWWVGxFwN5zD0MK1hMdsyDAwlPJe6u7m18P81o1zZ
MsgVyE8urEAPdfvQ1juerhs130M0AItUEWm2mlCQQxx25/LZvilPK/DWgjuTw0ed
sauCsL5TTsgCl7kYB7o8ON64Jme9ZQePk/AP4kkocvl1pOcTtdS/UkxjtiW/L5Vs
AYGUpsewQWnd6MlNvzVFPngS9yTZKbWGlrkb5rWUeQqgeaKxIPzwfLeGN5jEyhx7
zpBRExW2uCU0JhBIe0zfaBwmyEiPh1RAGq/WZQ3UAp8JBmJebwAcwMLNBt8BJvi/
p/+81aHlwJUF/e98F9b3sNzDAn8Ww5qiKAwH1H4TAqAwnPxilWXsNQ3Gbig74L4Y
hxhmmY85jOlV1ftJ3IUr8avWw+8kyvPVAror8oIHwFcOuQ0SyaIOGpj9H+WaU5QP
QJHdY1ZgGHKYoHrvfcBM5PQA8WT4NwJTSi7qhPJOCGez1BIyVafLxINZrSLt5jxJ
vYidpSJylSXl29wFHaVaDreURhtGe2P2o2CwPtGzsYwg8NFwTPLf/OEXW1iUieY8
ilCKPnuAuWMDctLvX3S8VpXmx/NE5gy6MXzd1NErs4meRp2YsU2NVhIdHNW3x1Nb
kmm5LsjUmOJA7fs3guXYw3u3XdVepMH6Mm1UgXFdnlmZQ/oClWtTm2TQsoY1KAgJ
hjNJ8DWFHPIysMPjFc57tvdXQCXDX/XXK3vzQCqmcAV+JPz+zpMA0z2JnVEdU63i
rCja7Jz2nBIEcMM0C3XVI76rW0TYG6NcyhngZIHeFstNGESrE57yqN3Z0Xo0eMHw
DpSWFh2B/VakQzgAwfTPQONpI1Xul00PvzLo07iIpmrScJkxmvTe6+pGeqENU2+G
tVSYArzrc3Y8x39Tu0dyQhHmqLo5J3KX1SGyR40vOsG4qsu28PtxR4DRXRhHwK4e
5Ilx3mSJohB9cNzPidoAWf38z/zfal+9EdfCuqJQTRihb0aQA94v+zVs3wWOhp8h
LWM+fzNmI5ugRLqjQCp+JjvaDgbbERoPGLjZI020mww3zohcJXvm7FbCklyFhAPc
vjZ/2ITeLrTa9yU26ohEwa/o9afzsHGAQb68AXDBY5Kxn8afBoNaJHBykJMPjiQS
4zQ28EkljmKY46FCDUP/4ummbDLfhgJ/Hrls7MhIqqfzUWFPMx8SdH+tavnYLEMk
vp52GzrODq/4YYZVPpO2QOzhwys8+92O+DCHsvvZx3Q6Eo349/nRoDw0IhzY9xvT
2EKa+gALiraHGRfTByok8Bszzg9ZQeMwec+xh+srwFSg4YQgT0KiP8zSdwMj+7tm
Ie4yVPsG1Eg3/kjVy0LR7KcS6uF/ADDYX0VUjTbwtA9KDc+Q2/MUMYa3FFnfBx5U
gvwKRLEgRDbo5L2s7HIPN/M2ueZRmHxNDJ1gEaAmbcFPfzk+TQ3T5PmMxzi0JGxR
5VrEuVu15okIFuCxRwWUc8KZclrp53UvJv/tZpifXeWmU/7IALc77m4oE54rm8PH
Rx1ozRhu5IQX/hi9k9yZ6/eZ6/mWxgeMcgm0ObWqqFu+iv7dVXi0tpZBLDP5k1+X
U1OOf/V91apP0yBllx+RJmvqhjW5LuLRDD9hk9MQBKsgGvXYJkQBBWr4YxnOPNL6
7XM3zBYkwz2r47oIyAJ7YYQcPdMKkU9zqAVMfgZeP4DfYjwjC5oO7hgmJAKKPUtK
EzSdDedETh/bzG+LPTWnq8fj43bqcSkoQHqD3Y7FFm9Ucq5c5DlkmjJxeSorPGnz
FLK3ZT5i139/8qYDJCo65GayOnItGT52B/INgsd56crGIjNIrWnxUvbxpjyty8yR
ONc/4dfE7qXOWyjpcBiJdcHeNj1hZhD2fWKfAQm86wN4VW7EllcK2pwexwAJNhCm
FspZ1IWwey82USxjRsLFcDdCUYgfsbw3Qn1WQcG2wScBGuz6N4s98M0q5wR5fn1F
Z+2EiPbwN92KX7IWVn+ngXl3lr/5xPa0cae5nJ/yFbUCEQivfTGxxkjoez1OB0nh
5qO5Hub3xTj3yrOwSge0Jn4vLl8CUIdQm2vXqS7AiZjL849cQtR/t41PxkG6DOer
ZEkitwCkrVfaVSeY1+a8acpjTwjkc7DTQTCSRiflsWt/yyfTrROUIoKnCc7MYdo7
bm1vy1o2y8Cd4h7absvqh+/kMtfXyGLarFsVgrmz+aj8zUF5LcehK1hassssu/M6
KECoprekTCoMl5l52APOkYiJ1F5xO8mX2m0GsIbba6s/Dfx4845W9fKR6O2fhBB0
wCq+S6iPkFCXKcJN2TaqB+NgFfIGX9ne+pCeyCOegPpD+Ls+eFXWhxMozRlQZguW
nbqqsSf/eMQlGakee966xwX1WXAh+vUwbAeRzfd0rBMIWk1b6ur9vL+iFD3G8W7/
oBrMWBumuRHdQ761t8VnQFI+t6SgNq0EeQZBEKRMuOL483t8XkoXGMzPF/M2OoX7
rL5MMC+BF0rlNrZb7HPBkOUa6h89wfj1NgWHhOAVoyZN962nZPW6JORdG/N7GIPD
482DlJ/Qp01WD5rEgWIEWSfqu44UtSyTbdl1N/aEUc0A5+YLhbxrTjxBIvUmyig/
d1/YjI0phvhrC2XyuvurNJZ7yJSpIZwQZmQfN4ljg9bM3K3N1anUmc2ntYTsQobM
AW1vDmwZ7UfaBRHFtSOiKn/wODQML+8TnAgHpgk3twQ1DOS/h3JPhv4vXXmqeoCP
8YBiwlVB2NzkIqI6gwzxy+OwwQOnPfcDIoRXTozYBIyUNiay5d6J2ZC1RyHJ1Ds/
G+DqJA+qruiu9MPMgPsVmyIap4AKd5IplpqjjkdRxl7Swz3FM09r5R04aFjy9D1j
jugRuDlP2ohdNI1nqqJufx7gfi6WrlpXZvMb+sjuxQjUf9wE2wlUGoT/4MVXSwPJ
pkbvhvSp9mlDNOzfUOYqdhb1/WSg4om+wLsDyBTCSOEhdqwN3xlPXH4DnSZKl8Ga
LR/r8jYe4CGmBZkCdBG0eYbKMs1UI1hW47l5oLV5znFGwFaMpTdJKPVwbWR3oih5
0Yt6zQXM1b+VY4fAaeJ6/3N/NDfu3AsGXTGIulZqbho/J1V4Pvv2Ha4jobpUyd/i
ROsxV9deDWwmhS806LwOO/xqphs1Myu9LtHYQdv8d5LFMW6AtGhXn3bZwdFpx6ZX
8KN8DzH6GU0LxtRRrBkzoCJIOqHV7B5E5jF7+q6vZcu5MbgKHStLKBbur83CHwUm
taStoGtKFyav3lMH8506S6wz6nIeW06a3L9rDLYLY/Bb0AYFsANS8aPBeKwIcjjI
bQo0R9QIabL/idKT4+yN0gSuQM/WtyZeKiY/AJuH2FFx47jP6Nuc4TlYAd4FGsFo
Xx1MTsVAI5lo/xOw4Ywg7wHQQiofs3ePB2KnU9m3czSc2+ZxzN91anyX28DlUTnb
fOBTKFE9EZ6oKp2WaCKLomjjVaxv7TMr2ol9eAXpNpZKiPUmftJssXDk7QXVdkYo
81eKak3yysK5zk7PUyx4uT/zq1F//9lDBdrd70LB6nFbC3CsseKbI6AZmRZER6Bx
9W9MkWjKs7wjhs4vnE3YRd8YY9QKtg+Kn9LzPysHtNDJ0ENOSNKXHKNSTjyDwWSP
fUgsVuXnZEP9Eb4FaHDwmxYePYBEQSSaKn2nprOUbQwKg3OHDWqQh+F5Z+TtUDSy
AqdU0VluBO3SFhetMieQJ30GsBewi2jsHqpZoR/Yrl70CSXUrhJ/nDakly2FleSC
OEySK1H6cBoH+RpPHzIgONQcz0lUrjOCB/CSeto7iu+x6CPqxTk0zgQLObp+IeDT
D+ByfMXNNn0E1Q9iSJVIRqUh+7NnTKyljzj3Ow84q/IxTZLrN6YUVYlYTPTUv7Cc
gT2KMZ/L7DR5HopsJHgvAv2SB/BehvWxXWBiW6oUEp5RY0aKd411/fQQSuHEfOvw
7KCN98610yAb5gpILik0ssy9YhOVZGWcipyE6nouk0jIKVz6HwyR+GtS4pS2lYnZ
nWXZb+OkuMOWaqGWGEaH970LIt64zzxOuqnivxyfHxOgJvV6FjtFQIAunHuPA3m4
vVkDAjd5fa7CIyxAb08eWskUf6iwivowGzuPQRhHI3FRw3zL22sBrkuILumpapLh
fwOWPSntTNmAh8Nwg3AlV6zUAOlccbjE+zEmRpGWL0y6/iaVGLMeR7F0npwS7Tro
lUo+ti1zzt/UBFclM4xlNFQqo6NuqIgSFwD3k7p76JrzJkqCJEzxWHMiO/nZ8E97
HEaZLg+gw5Vahq0gdQ9g0AUdkzGXNXxw03CbVuYtTLFDNv0rEP7/V3ts/N9g2inT
xEr6SydHloEHBrxb8zVBP6EwhIlq+ipVoJLEkuYL4gU2INnP+v/slZcVQOjsbrw4
7I9ij0p+5sQmZmCCrqfOePzX7lyEbNegD5FpB1p3EBEWL6b5Z8FcsRbSxTYDjvU1
vGXb3cVM0jobpzSgPOlbr6uXVr6mcfeQtKKETCdoXHHdziflOpmDgu44UJBGzGt9
fW7SzYYOIUec98w28cbSJArgLFVLUeWpLcYudrOvyDV/5kHS1gdyppmUzu80Z+MC
kv47Q7WyRYCHKJiP+VGX0fNbqvLkitn3EA2cIk2AHO2wG5KTzhllzFtV72TFaT2A
lAHRt6/0VybHXumZk9mxPhbeM9wNR/cbOWyZp16Ro+hBaenYsVtWFw/PYboYU7lH
xdqEwK0ukYfsw3XtNiiMYak8brXAJLlYd3dpIWhuD1KIff932/9+NaCarEQQqZvj
x8W6FY8MB9SNcX88tarIKanp/H2q5vmNbUam82oo5w3tqc3l3ER0L9TkiNGkYjP1
5SJSvUR+XTmG/BIAZ0YnkdYttZqIKQWamkDeZNkjcNFZynvVfKw1m2ZeM7sc59S+
gjYMcY5TqOBzB6RSGomR7qNB2Phj9guHH8nY2sBVsRY1UxxrX4+yXIc0uX9LcCv4
bAXHeHhes7PJUDFAbJE1SwlqMpLpOkA/TsbZ6zAXAgKsyfeX7YSUgOjCmA/B3Nwh
QLrKlh9QZ19aXHfvJTxq71CWOHR9/01vpDrvocgzDin/WPCdZTOtXIiYJ0RdnhHm
mQpFpFkLL9B7tZ6iprTqM5bFpC79F4xihfxURA/vkI5SLFp7EfNUxv5yXJ3PDtL3
n1W1GrbjZPd50jSch3tkQISbtUWzfD4GmgzXhMW8ycviByF3jVo7/6Jmj+D9vCBw
g5tmXNKdJ7uceOouiSf/FgPmrJKMZ/B+RmYY1m67wXEezL+yBHkdv9BzM7CTJ0OL
7endWr5QBvBwpmw535w+WdkSurFlaJpSYy5uW2xNF8RN7t+3gHZs0PhayPCPnxVu
d7zJOgPAyvvy5VaLHS30eljLGheUi3412mquq86XA5Td6FpdaqfboAhzsczT9s+5
579JfscQV2Ok8w1yX6R35ybZTx+AF43oLEj1hVJRS36Q6DQNJJECK/50MPHoipKU
WAUf1Ga5cBNLrkuGwm5G51JHub1cCfzhQWDfUDRuO3StqDmyT1RGt0lFugYIE+E8
RQrvEN6JYm5c/LWFq8IWuocowiv+IdMZ2ZfpIn7bqFjc40B3y/2G0Bb3eKhgORwA
+7kbb7gp9VlrUmvP+q9Wk10qyylQE7MWN4NY3qibrgXi9+ABISkmqbV7mj/wZrFV
616UBEopiInifVsuQIWbgP1iGDvfSaS7qUHNZ7dP+7OnOSI2my6sq0c3kET5WLf3
t0HZcN/VkCq0o+TXQ7Ck9ycOn1eHXIJmTslBI5lr6dj2kchII62K8Iri06k32FXT
uKPaqEohIQxsF0IRaglNlM9FnTYDPecQlkvx1E2OciJz1RAfRu2ozpAwCQWUWQFZ
JaEDArAPhBSlU+1jA9uWmAz3w+1DTnqvqwCKwbEd8Kx8nC/IWMfw7DNEp7enXDPe
l5ic3NVtZxzJ5z/X7vD+5HV3kdvKyf5muWufwyaYmjo8bA75D3PKGGWjMdwUlow2
jm0L63Ub/wlHWAv9yklk0aB39qBxbVg8+jZJrM0ZMlNITZVxA5EWgpilw3IcBjCd
F8J/XVEQG3I/K4hvGDJCx7fyYFEqeQw2hGTaR/cYkb9Za/DwXtLbmXdAZGXNySrC
6fNy1TJC3kikLyyDba3B30rbezU/ogmfSbaa82bUAJBTQLj2raZz0Ba53AnYr3JK
bDioQ2Pw7T5EW29t2s+l1V+O8xBgmsAOR5FH5G4TPmUBwK3a/Vd2CZNJcWjnTk2R
0iqULr1tJ1nBZM8fCMhQRs1lC/8IksrE8rzSunP2tvk0OyXLaKE3bBflABLGBN5i
qvgorU5sOeW4H8xK+CzRrxn4288CC1f7V97zmcrV1I0DFBjsiapuklgQ+g28veOs
Yysym/Tqh5AN8/S7O0yclVKDW1jFlhAWlA07zX0U4DzukDWHBfqjqbvTcYgToCLb
BRoKpCc/ehFclgUiDa6WU+nVjiinaIzLeAG4vX/YaPwA8Y1rrcZmdgPW+Z3nS5CD
GzwZKAPeHZ4B9Z2dEmba07SolDz0uuafhbb8/IUExvw+nnj60HbLPO4tqCOohGlG
tj5KMjCNImspukBuAIEO7tjMZab6HF5DSqf4Exj5sETuVW182UTXo9oYETyTUq9B
Vjzy5X7+T3ZrEs3r0Q4E9CdTDLu5bc2V1Y6NgtgVyi1eQD64iR39+bV3FkMWX5Yy
CpNRKnXELhQTTmTx+YKiLJooaGrMVfhfwqkb715O3P1laG+811xrvB8Ms55Xy7bI
KuK+b8CuRDQlUSXy/Lbj/u6JzlKRQ80qds8giFgxUJJqwsWUDu67EveX8bXo188f
NAcnGf9egODUp5zq0bBG0jjruiDn8vhj2TgK1S2R6/hcfZ/tPmpMTGsEAQ8BoqR6
20QK/sBPg3Izc1WjW67EGqBCz6SXsKnwIFFmK4MnaOwB1WMY/KXtNJIA9twgc2Jv
GixoT0/5htCFkqVuQdwdHjtM9JttslhVNa7dato+h3BVzoRIUp8C8d1g/6wx4uqQ
ddhODSBMJutYhVypLZj6Wvnm0ctIOnegqsqr8t/2II8/A+P54sdx+Fhb1GT1LEWL
Ae34qcSa0eBwxsxcvc8b+RYipxJ7L8m9EhGZG798Xa3ZRKn3tJRYk4o1ghit5Sl6
HjSKoD//4gxR37zEkyuQWAVfP/jgko7fIhY5ZxK+TQ3pa8srQmUZJuu0PAWwXHok
gMTmv6TN7ia2mziBLAKUFGIpRcfxE1IE7QgBPA58n9NonDsBA2wZUvWy9h4DMmqf
odpXIA/raUEifJoPA5kVddaY/0vP3dEasTt1dMnAMHWdRpNpz94GMVGQE32J2ZwE
NH4rpOw+5ksjDDt9HNk0/eOM5fBXwG3yhn6CeUxGlq7orQXenXxpf6zllIzvD3Vc
zkgDF4s8sJwXPT870fXeSOH6e54QvLy9LS26waR8uoTtKa5BTmiILZHy92vmewW1
GXmaNG53YXL4aV/8QUMs3WFPCsyrXrGGxvpMqlJ89B0B8NGKkaLSWWs00D8Bc9j3
qPus3BBZX4IePvwFNjE6OFaCGkbM4sJ4r5Lh9FFVHHP9xDa9aVQtOP0YChEiqapi
HZdhszFwY//NTd5mYaqR33X1k3zSE7ad/xCKtxeZoUq8InK2cb7F5D1oDqou7prb
LXhf2VR5s9ZHi8Vh0k78BEvcW3obKBxZttNinb00/Z7vwBfvcco+KTcrZ+ZznF4V
C+WVug2OWsJ4MrGVS6zYmg+LelLpOzIOfLZ+tgji0BbGDhNIJ5zRG+QcIUStduRU
Kn63/PGctnE7pSZZFj/SLLiPEUq3GEBTXaSPOT1FY4N7+pkkcuo+KL5dHVRIlh+0
g4DDstDfHQ9s5L0wINe1nkUqmiC6ltyaG0npVL3xZF7fwFqRB8fCDJGsd5rU6bdD
Na2QdOwidKHuUY+VCwmC5VVUAJR8LCEvhBjl2U4yJq1Lzm6JB9Bsmv3wki2VvKxf
My3oEYhqpx2Uxn4X0DyO+kNZ895L6k181zwPaF0s3oNbQ/w3P+Vcqm87VMraroIH
SLCbkyat3i7wwCeM5/mVBay14tRtIpDH3dD/XF5rpEmyjI+12XJKqJIIJDDS8Izj
Cbe9kk5KgxrNR3Fh383xJxjTN9NQVY71mRd0OkZn7RpsGx6tbfXdtWJ34ASkcReF
eTLcVXPzvRIILvq3EORj6wKlKZQkUMuz6M4XDgs0CTzVW3V5ph1xfWFi+JY3aERe
AAFYLbxUx3zDc19I9vd7m2j4Mc33C3JM9JC2MlRQmMEC/CVHIrGci/LXEzjgEqpg
2lqxTpO9aryFhyLAgy5VLAgXMzudB+H0y5sOITuO6TFkwrQxItrE8IiyTWy2gQ+w
7LIdCfmz9byiQNoiSIjxM8lGyWFtH9yXQFAqW1AO1rINDs5dqNpGSQ78cG0KleFd
bVxUQT7C4xReP2A80aXQ6uZwLv7e1KSzRAWy8LdZauXNQAl4eklsjvyAv5BO1WMG
/u/++yl2iez2bJ5A40n503tJaWVQxxKGyWo7yxyvh2K1mkgbrWtOfwSH4AkzE83H
zZDHjubTHa9F2whHhIFjVRH3jWseAzAZxUalfumy5+NCnA63oHpU656VPATjXyG9
lPL8gtNTjskc1omJf1Bizrjv3iCeJn4CVIA7fWdWc6kcugK1mwXhmZrn4gzPeRLE
Y1MW/OMiCViWv4TdXoN5aGa44cdAdr2vmvo8K5zl4xI7WmPTHarAm0yrOksJ2DIe
m5eZ9DqJQJvJOSHYumpl4INEuXhX4NleykBIdqhobG4fAlsXqCdtx8Hn3wUkZuVf
utM+RTQrhJLgZYca225XUrC/MQjJJkKEI+Q8DeF9VBeNVC/wGzlOxUNYqYz82EHF
fyWqjHxbZjkvoYtO1XszHelcJv7u3VCcXyue4gYvKVe1fZKvzCA+P3FNV3y6UDmM
C2JIAVfcwR4Egp4CfspcvYW4hGz/wFi2Tch8+3PEo8MhwxlxJe1R1j7lzmU+roPJ
MTxgsNKYuj+BppokQtQ7DFEecCdY2USFaCL6fAu01Mvnd0Xo5RwBiCdPZ38zw0T9
ubCxHG9T5G9U+cVdwnvZC2YRC5EzkMJe5PR+2IOIL/3gsjXGRifFeSmxTLnQehmB
H+fIa4/V1IGi/4ZN5/wq9tw1kBVlqhzi98inUDVG0zU2dtwnMR9YhoKkGyO/mGYb
/xd7NRbHCbR2JmLp8idPu0JCAQxNuHa5yE8rEK5f/2FyoXHGz1nIIH5WPRIADVb+
0DigGw/G2T/5zokfjhim0Hgms80f2HwABWfP9hCz6mBlheJzs0IEVwgrkk0en/yb
qsqdSgxxpBfkkRo5ggK3gA7Dfsy8s9NV0DUlAQPLtVttZuWn/dcMmdUBWvvTNeyP
nx/WfzRnlGAeZ2v7GdYFtXDKdHmNh4tykQZeNaXlud9E85gZy8nnrJHPm0iiiZXA
2gusP1wAxI1JpnKyW0D+IzSAuU057IwxWL3lnJs9+C/g6oI2XqRPnkkBMfj/uL/4
cPno0ElpFObwqqB3Utl9XmC5KmfrBzYVDOHxhOyK/Mc+diyqyz/9HGL8kJ6h7Ldz
dwSPJOEFRs13rJVoEcntG4AauZ4tkpeXVWe/X557yuk+vWaY7MPiXJG2DqXP9FiC
jkUsD5Rau9LCiYkChIm3OcokEnyy10PVPtbcWud3wSsQkbSgvcB4A4uZ4LnWd9I1
kTn0EQbQqKkQw0Gv5gvX+vVm0/X2H6LTNTNB1utAn3bhxStAV2GvCMHwTbObbF/V
9U5RubyJtzjOfpRBiFBSfDwUMDfRSqShgfE98TtLbhRoI2k2RfyOFd8T+oeR/gfe
cKaFnu9dVwVvP/SHlNblUamyclcKhwbAZdE+Z9WgNE/tgJsOSP2majGtuugOz9fe
DKU8Lj8NDB7GTlY943sQ1kzhk5htEfAcMjeUzW8H1kVgmXOWqslubE8SSq3xZ5xs
InTtJNS67oDZnUwmikuy65BC8vfCf8nqK/062gyvZzIYOlEHZLUXUYp6O3zYcUBj
k3oFdRNsH87e/kHlDN4uUMDsU20RisXxli8jWvtZyXrlOhAp5BgF4n7bnfto/XAh
IxufC3eoxSQWQ1VuRAT2+qR+eld4Fl+r6ZNMoDBci1dHBxyVgnL4UeVzC9XtMYSk
r3HAVJ/5uS3tRad4tPicDtSf9Yix39T7J1mpnzjuYlULvViI9egMAlgxC7I1OYFt
qWAxgnkw8EkkOtW4ztrvqluc1r5PPuU7GinYKQSuSc9HxM95pfEFawvWJNqrAP3X
+51mqSHIT5ifcxccx1ESww+Kk0HBrIGriRLYXz5CKz+s53giSsV29MXaVLaNiyc5
3krF6BJwSBVEprfbbv7tesaemh7eCMH3nuzu7yZ+5FS3Uuslqp9rHw+oLp8H3TzF
gGSZLVBGqn89fdwkav4ozBUu2EEF3oWiSAtg+N+mjYwA5HHg+3hjzwqnw2rIEELU
K9IWooC9M6TE3G7WoasC79JkdEMLnB0CcB68AWeHmyR+Ko9bcTMDn93l6G+Q2uiz
FuQfzzQmqOZ36+MJF/AquNN6S7AaPWj1FtzMbj8mTFuM21mJacpf3SOEB221GyCh
WTCHQYZPAZEhJhJWfFtuq5pqZz4frPZ3ZHPS0/VxqDxpk03na7z0gouEStOnVFt2
4WfvojrR1lXsvfXTOLe7RsxHk59jV6w2cYHjPOr1PMd+5u5yNIvoZkxLJ0C2G4TW
oAfoWeZsnlvSztRfAGgt+bXrh/KqcMJ2Ag1ByMNTmx9tdKhDdKaGkXCv7mwahbrI
Vz9/qO6qKc3YOrwi5/fjdF55XBFwtQfdJ4alI+pQhXLGlm80DTIM6Ao6pNVsErjy
AsmENk9b485WwG6I5/54XnAq+RLWI9kBXwt9/qbxOQwED4UMKsMKDzbH+oNzxTXu
RPhUDYtZ+yuo1g8DiMfSbMeN9EON5TzbR+it8q0wt8VzhS/5uvbMQCubg1dpBVMp
VhlttfDY+7S7H7BvWw6fcMNN5Y4zbhmfD8B6dl4OlDiqA88GcPDE0u4RRY0PxZNc
m+4h3adCgcDftWGC3na4ggVZTAHFewWtL9PmEZHaGA2C0WRx5supmj1d4TRgwQfQ
t7YSGScWNFaMxUhBi5RD6JsjQLmkbnaV7C4DHx01SFHwYffXFzAk+wjX6gHyOjkl
8UrlmBA+jpcWgt4fAzqf/fk9Zy7YkWjsy1vVmkTqT4sp2LPr4g/RPuo1wn4Aa/1L
IuOxtXSO/T8CrsGAGctfHJp6GHCtyZ2w4cYQ8rWxhKOediyLm1EfCguadScEW58N
mLiC8H2L4JSp84NcB2CdM7+1dLLsijiY4NH94Id93bJs/QDrYFzceoM7xCIIUxLw
jf8xCN5hIPdctByKuk64jeXrHUKhAO61uPRp+2mtfIIx05QlTwod+bMHz3yqYXdV
aONi3+PYB9bvacBmvjL7IxJmX+QKH0IyhEIMqw9oN3MFlFoHhwfAcf50u3sMnbps
Ytmi4XivWEB0jC7otIPVmv1KRB8iFwKpcA4i2z4nIdS7VAqRR7GRtoD60H/Oxlf2
ce7YLj9ZDkLja4r6CRBZQszgXQNR7tjBvNfRXiPsmJbkAsUfMfwgk5zkgVRE6pcn
4SisKOy8XGFjHorGHdQnUgVczrpcdQvSp5zkn0zBsSFPYDM3OgBE0aNi5NBxujaU
fh6HYkxuP2/be15Y7LElUxoqSduE+kP5O3N8VXUBdB1IQT4cUooaVfUt04k15xU5
/eilX4OxC3UFLp0v6GdVnYAKLomFpXOkteubhxzGGs8dzl1uheahuhbD8xBZyMIx
gLXb0XcOIDThMToiKU+PYKaigSFtKFysNojGT2kooHXcia1pJgq8cwHoCupc9pyB
dPJODt7hMvnVAq56YaxtRd2LzF4jcHE2hZRXesb/Qx6r1seSp5nSmeeP8EPbKCA4
ZnewuYrASXCsf4pfyiam0X9bhSQ/XBNV2zX6ll4zYVsUiPYQpAZfDjcu4xY5pHlB
sdYvZG3p61uQx3IHSV8dRaB20hmICe7VSsTIZYpNm88pYUsome2caSforIyStXQ+
nw0oT98gAAzAjF4HGcv+rSIAGNu3wZgEtAr5tWRKrC48iUmypUY05fD8bHILLGso
qj+LlmAFnFPewqfR8LitOnj0nobWpwZGH0zW1xCAVdp6B7CP3un/GHyKfDfnz33C
EX2LqVy3rWyZCrNl7SWvgUFqAy7GTiD+OxewI9oTWGXVnOkvRECr/ANFRhdrXifn
w5O4TczMuKkOKWQ8nXwxUikCckliDUIy8U46TLNfcKNX1G292zVMFOw00fMwuf/r
N92Cxv99mXGTuySa6KXqWbI33XJQ4oAUM2QkhN1bPvUNHWTLIHPmIt7icn8hWyTJ
44+k2P2M7yys7id70rRchEiWgIQ/SdqTiV/p9naaPlkuP0uAX1CCoay5qZKTTXv4
Xy1xskUrBaVh6zQxx/24cfaypkhN7Yjy6jnQl4Hf5ugpegvBkFMzw6oL5Y9Bi8yj
n0aJeVSqRJKMWjmEkyFaSOB8wYXFJmNR2ZsKqFowD7PknumLeRStafUORH/KCUtP
nLPyYZj9WdfZoKZnfO1CI1zOtq66PfTCUXGLJNL0MRpQdSg6vmzw9alFxmGHWbDk
VGnZYEjKD4ULO67N6JPE1hzUfWkErDZgYDEwrqm2kJsaa3Zw2K+/BozzIdQrS4M4
/pgvUA4I6SyQ14DZe+fp5xKwPf2RsRXsox+0oO8wI+Nme8QiZ6emsUhKmsZwDfdP
n2HLcRTNAgqTzMG/xZTUv8k4kpFSFpcVDP5HcKMhvFIqlXDYatL1AXnsd75elG6W
1fz8YkYVkNe7Dfm4d5Vq/Ow+8Olp5QYguB05oiqIdgWL27QV5vw/BsnRp+FbeKim
iHjwR/xt/m5LrBeCoEuonMvrC/cJW+GCZeq8mIC/NnCakcpNYDB+SEPJJCVjndRm
BcE3tY68WZrRG77TxS70U1rfObZ5HUU0FNbmX5MTWd3sPM7blnKGQbnUPAOUaBkT
JTpH7G2KTzkzVFWOT8nsBn1jcGhULQ9lJ7g/CrCnYCYBH1kPfAxkMCQCUx2b9WkX
GtwEqw8oOEkdhh5uLKlFJCgr+5izYnXexPelIZa34EP1NvCOIyUdVLKTKP8YYlOj
qAd3iIK8P6PpPJ4WTayDUJpxrLWFGo0pegwZk8oB1pxzfRZSY+iOcX2trSyg0VcE
QZR7VzWc6BROaJxBqbAeqh/cmP+fqUH5kkuq87snAeLKcioWp5/YWL+gKLnOJIM3
lMzDsqw4RQ/u3vpT2COweAXhv7GIrHPGCqHM12INOF5mKvZ0lXloyFZp5EwrNz/a
amsCNuqzUgUkiASSAgsV0mHKIZnxsHp3GS2JuzYcM46J8s1XJCrRnvqhXKefzByk
C0IPD/p+TUSSZ9qzjdDnUFwzGXUfsMRlIEC2iB4YuGPA7nFS+VBHJZ614reCCb9k
+Md7TV8G+ApBwoVTZ3x/saj0RqPz2DJQUnrXHFF9pI5GCZtKMtmupp9jAbfVxRAZ
1LgWa6shQ7jCuhOcVeSH4Yc4keNSkMEIoYTQiWfPYjLzFVVGmEb8M8v9v8xMKK4h
kJ34QPFSz85RPbliM/AX7gb+7LgoETlykDJQLY4VIt+U9KLMzbIo8/TBD+zGtq7a
cuiA1pcwzjl8rqqseeqdCTyexXhG+pBLQgLQ53QP21BNoKD8WfUnw8ExKHp+zm5p
2JJicpIG5ZA+2zS/g3HIVzF3A+S0MKYZE9ExeiJ4YfZJBz9MtQlPiBa9tdPexFYo
tCc/NQZwdRfZGpBxg7jBhGQpXCJ2GD5LMIhWk+gaGlOxx6i6u4hJvobsbFnvrtg+
7ueM/uc7e2tnPgmrLsZbnxD+KkLXJcsdn66zbWgBV7TBwG035pLycCanqGBJ+xUc
vFKLAN8k/D9nuwK5kd6RleBGrQaGZmYJBEsDrL+n8eejZGGUbj+z8g0S6AlAJJeS
vFNd/6ydYMUka1nlRmNTtgaD5xlAEp6dU2jCK9A9y1oD6l1oKcFVAxeiOspPifLl
812LpJzThvSSM7E24VyGRKKOWMb1TMpPOTFMU7x+xO6Wo0JmrBBHw+Cy+GobqN4a
GSiYZ1O+7gwixy4oud5DdqvP1f66maglkPLKR6K+nYMP8di34ljXfNj+uhVbI0KV
8H1yiVK9TQ8mU4tjcyurILucCDgO+znPFZbM4LUU5Kf4K/sZGEGOOWH9m2XsWhT8
R+bEHLblaOGCuWWEKrmsHej2ktee8ld76QnPNKc5EsVgCUk1sXcDOn5L+G9sIyfa
OOTfnu4Xq9fWJgPHmx8n23N/uNYYWwPtTl/uRb0rN5uBmM+zLh3X/XcfGtlkJ1IH
rH075lF0G4R6XqnufNTCrP6pTcmk5u3/V5r8N9NgIhUOCRG0Yllyt6gnigGaOixC
kYcNmX80yNOybgzFrm2BBq3riTaO0v9RBsUPISuK48d03xprJjN6Z6JxpEaoNj+5
dT60TniLHaJ7NdtsMTBDW6cx1Vi1spiSXbimSq4llWqpqYbmdCnP8zRnFc9ww6M+
FtEjyYnmOow1hhxhcvbNye1V4h6jPBH5DvHjhLh2yUjwmsr7sKbE75CHR3ejnGCt
1JuB/kFbu2ktuGcxVsk/r+Fhayq+9nHPuEAV22N6CHPaE3EX46oJ/1anAECp6eVu
6C/VovO68PqcsBE0fYauZ0+TzP8wlLLJazzYl0nzhJQsa45wyiIqpZaDnEpmlDkG
gtYfF/3G0qCY0HN4OL6e0CYTQdeVAQs9cm4iOHBtyMSTrb4NZpcLRFpo3Uj8dCRt
Zt/hGdaqQm9djsU4ikBd8x7f7VLj8ue+iNxXAki34b4/9n/ZB8DlOLZwz9GIKA1/
g7571FktSU2h4Ve78hj4vdw39FbI8PnhJqNYpHBmFK3Pswa9XjOEriPpx41ZC/f8
1CwbsjRogWY0kYHNLi/bUSc1U58JyUu5MH6eX5sqf23oj0q4TBvnk80ZaVn8hOMn
qh3l3hbmHUEQglRkKfsgrpz1/pdl8EN8N4zOCHCgcx5T0fTm9ISOH4eAHhn/ssiQ
Kgb3TQfnGWk3E2X7EF4zsCMVgOVvWYfVdqka5D3VkHYQ/a6iYgoCVzPD+zl6eHz3
mFjAn2SGi0VSrJQmIvrvqeSgWfIxjsr/Bwp46UnPl6VNnchwBB0w5YxV63S0yhwy
eQl86uMb3Roq895VNOEF/MrmX4CERzE9hfAI0unUXnAEGZlaV+6ipRdXhWDIGK6J
v/yhoCYHoRXIIe4qRigjATGFCUZNIG7DI6M1xWuLTHeQGowwSwkxgNC90EzcJolf
txzx6FrcC9lmfHj8mSnUwdWnxYdUs1NJyBZNnMALFJDveOQ3+bncProj7pg0gOdU
QRM0lFU1v+o/Qfg28PVGuWHOn/p2yQPS2HC4zJ8klYh1vII/fdAlyva0RpWW7NRH
vemGWuL7CwJV7y+HYZzbyln3eUdwb7Me/YfxuYVJ/BlSMz4lv+mOupN2IJjpE2Y/
QNOPwx5Ne9CQfpPRuzO3MPNuSM2Ahe45XsYvxlgH3nNCj07OcWi/2MtogQuouSzW
nFaFJNTpCGmcuJqi+BADUDdDbB10lTglrAfBLS03MNMsei9wNxsW9Qu/jR+RacQn
G0XIrqWOEcQOpX4Cs8r5KvNoigUvTGl0P41TbL121ELN/lAYWkGBcJ2Kpp1XW48L
rWYfR12w9pjS32BWjXrKUVdZUbzMIwbuJoGV/0fnQ6skY5Gd2CaT9Wk6SpP8XLKo
Rc8IvpRunCPxb9SxIdzg7dg44vbi1VQOky467e4pGiKOoQM/DZoQHI4HeQOyC/Mz
4XIlZ3IwJb9MU6E3aUJPp8Sj7ILcdnyfhxrGXB2zTF6GN6hbsmpB1zPIZ5bF/A3g
U6FAGcQL9aD6aeWTSmOmLRS1su8YrvdH6qMqK7hAane/fPdMix0sofnnYe0X+Gcr
R5C+IKdEZcoEV2AMiPPjC2r4RmUcJwnVhSa263sV21Ow94tSRuUjzVJLEtAnGADq
ptZFhWsk1jH4IAMMJG+eJRExgUGaIyZ6JrVvmDZXwLGDtGB0Cf61B6xxiG+o0uUB
b3I1gh0mL0sJhzGLHGq/dJwV7QUQcBWVEg5arQn9QHk8zb790wTVv0hT0184Btr8
MB//hng0L4xa38yX1KJM/Z0eVzs/ewqK7GySJ1nJw6RVCyYFa75eScSnYNnuQMAV
ZF0lwgAz6uDIj9RphhEJnjbq9dUaATZgAJy48OYhc4PLseF+7nb7bEroHDg/gB3G
cIOcjVF9663yfh1yIRw7N+X/yGkxhwl8MdjQF/CQb/6wNy2YP3LCFkmbtcqL1bte
ArBx60mkaUg5OfaAJOnH1SkeI7Zjx4Qw/taqve+bhWd2tZiicID3EEPN0gSZrMnV
gsnvRzxlhlZK5Z+QS+BiNBA0HtnQ2jb4HjcOjNoYBoxQFSJM3fo4DS+rtoNIPcGm
OtJHuy/+CfYumX1KH4aNwTcpztMdac7hupWVqJS+kk1yCPZPKI9uwOsP++IJufRG
g0hpBPihIpOOu641Zc9TbtR9IMtW+zfZYwzLdBB6/a06bBb1gQMUUXEjccxIOWN/
bzS0ZFf/BWu3qZAA1a4BiE8fEqp4Tw9onGJ6lgtT/ASqm8FCa11ABr1h/NONeJsR
EUwGQwCV8BneryIxufbZWPiNHjtx41yDyJtUuwgywYM7OAwFQYBQeOQaMMzGMk33
OBE82xqpOAfgpO8YaKHqKqKJG1ZN38PXR1UzyFPuN8zkLtDrdFwxpgrbuN76qQgK
O+7pHcFJN4EVaf//E/7hf/+Zbueh2Z7dOtfhenmEcNwtF2LdyizRetojdgXHuQCa
BKt+IlJG+ULrGTqii0qHgKGJcnotVj3N8eQhT0C3uM5uBVA1U+rfLKqkzK9+GuP9
Lc9U0y8YUrMdZCYO+J2Cebeaql//c+V2S5O5lykWxRNF00pL5g8sAve41uj5pfNf
yEOukO3G84c5JFQjtkPfT5flJVMw6laOAbPpvw0fH5u0zxq3OyXt0vzPZ4vVd8Wm
hYItz6DAfRgssmfWzNeOy1uvBRbQhxHLtxO+Lc68OVx1zTko7GLJEuQb2nW6kTZA
5ipkaq2IRnXXCFvH16g5zIU6lgd33rzDhBZuVHJsSKjp22miwuC/edtdLYRCP1F0
D/NzYGXtEKjuxa9o8ju3h22YXJjh0AGMOJPyzJPw5nibrbdlvP8g/s2g0C/VI+VU
c+dJUK+KNGd2wXneStgEsAfhkKyc1JvkwfDOSArRParxJcCF1815fRtF18YurzIG
8WdFveOXbT0NgAWLebYSUfdIaqCJusAQCOlvCb3wss64cTLi6pzcLgJEBRBk8xGN
68ez6H4rC2F072WXneTrwxt2dWJ+dqnfsEQb3MgaHqis4j/GDhNd0oYCcJPagITd
ReEskBBg1AK1N5Xc/DrIbgHOEF41vLMviyEugkNX3J4CTJdL7JLBbjGc7Z43AsGs
stNo6Iln7Q/IL0zuiy0iDIU1q2agGN9qTUryPw641XtG+QWjsTqb1MSpJR98DeWw
1YgGSr039MEGKco4sEbLDvmKS5SEUpBTdnSYZFxArVQZoQCbtCpe8JuHvrZuT0al
66BIBjARAx/kmfDR7RlxY4oHCKDla1trxbWgG09NreO38Ho4FTtvDW0KGB7AaSAF
l5hdQ4d/5oAWMPQX2ZNqGGfoKfoV5itl3bGN7lLiEhQEnEI7BOitSeUvv10wyUIV
vFsXRvVdWJnAg0etbRSPl7wdkV4cnrY/9M/8aiX52fMRcKvZx2FIU3/xP5MMtg5n
fP/vIDapC8Wqr6OgDYsTk2BNQNOIrWaqcRtr00ApQ07GVg33ooFhOl6CYwM1dlh7
U8bdqn2Uj4b0YDXaJVcd99BJTi7lCdzUckggcQufJYm6RuuXFokoV40iUGyb0Rhx
oo3rpVVBSUhO57pPp0qkrSreKEB5KI050H/iiC7R38NaG+fyy/P+B6sy2WEY8niQ
XrsbbXhOIBG2QJmSMsRLHL/Qnhx0kEMj8h/5loIdXzGfs70hWkRrkVhoUr1PkJFG
PVAsbpbm5YZQ37aqZGMCaycGv6UAqnNPJyO0bb7bQz9WeMwt0mJ5HaLrRHG9Oapm
H5fwaBV2vVnLu1B1QaQvzMZVrFVBwEofAuorhWhhcZvrLt58xiAPWPitEMmjVK84
iPabkJ3gDRZk+5lF/TN5vloYRrCJuEZ94hYV6UEE3IFEFV3TTS7UTOjYr65+FJaK
Wxma/5cWc6J2v5nsoxXO9CnGroqs7RM+cBbYLa0tsWHEB+SWOfkW87ypMYZYkQ0e
zzV3ry2kR+XRLqDJ95fv6KTbb1K/F69BsWMNbexHdSllLVKQsHumXAs8J1f2WULV
tqI61dZ0KVTgWaKwGEnzXNx/lJCvkVuccgm8abkcKOBtyuR7BXdkSPWZVdnt3tjv
bqDruMPAFyq84U5kNHtZHDIdCNb9Zn4Ks3Phkdyr9cuBxb7TgDGoaSZ3yHtBkBx7
dmsMw8BszbecEG6+PkDBbt7+DJweh55knOUDVqfbVBBFhxw8WVY0FZx1iIRtyFyw
xLtB90t2gzsrYWbUCixA7E/HgoBm9Ao87nSOU7GpVbLJNFXTDPuK0QM0Dkty94rz
OhkSbfdZw2JlRFG1RA8ew1asayQEbWFc2P7HifL0zPHZZGo9aMVs5ZMcbBaVOp6+
bJmaT176p6zDLiMZP7v+jCvXyh5u/p71EZjrZ971y46T3hL6x+AW85+ceFSi3ML9
aTg/0XhXBeE5rPit3tnbXh1ThDyqI80CQa4zPuW1hvdnPLLkIuVxaXObsSJCie+1
/0M8ZLfYgYFy3Ij4gPttGwkUds0vnKmGZUCeLTvhNS03NI46hG1pDentaWaSf8vq
dBgBFtu1MYrv1kI9LUmw6eeIEUEf0n6rSgeBCnK2QpJDRyxL+EF6lAx8I01739na
cR5ZG/RXw5tJW152q3YWwGQQcLGy2vsicQ6lkX2OE9PVXQzuUQgW9uuWxD7Io7SE
QMbBbypnAd8ueS4QrWL42TFiGd3+HJMDwQWbqKcjZuivyXU/VHjsbX7GoIn9+aQ8
DS2wssKQmbQ/Q70bEM7lA/rHY0f+8HsX+80nMw+H900DA7drN1R4UqfGFvIh8Tyh
HLCjq0S1csfzGahNbtin0ZNVrtuu33SQKXBXY5YjQeoeiSu+60R8QEuUUbyYwJha
61s0knjR/zzpu+0TShyEFpjcE5roMH78Hn5ZrfioyJmNc8xKGRQjvI8kHbEnJJ8c
gBhiKDmbqbxJKKUww7zR7nI0WDtJc+WrRb78PgLMmL9UrZWiaCkRfptz9FTNC1Yg
YAeJBF840omTTFTtdwh0qovWIyjOkhHnEvomonjItOdojFsaXfq/u2+F/JMImMs2
MrAgZg+LytDxnD2frmgtG/0ODTpnkqTj7awW3jBHnxJLKe7bW3gftkSL30TKjgzt
fwunSPwMdd/O5ZbBnytLnE/qP2X57UyXiskOALk8pUJlaXlFy8JqpgbB+7sJ2EcG
mNnt3c8YJkdkSFU/TbHFQPNGMbOuEsNZlAnPA2B/c+Qd6jwGd4NrNvc/Uhc1aHEp
Khvpi9Lr5lG1djTbg80m/SOBfCw2xtCjH6JFDkjCc861kXzWMIpPVT++QTsYRh2Y
QJ4uDyKw9+se4OidGZLCMoSP47sow/9ckU4aR9Xztlkf/HupzjSv8PyAUWOjjLQF
DphfuFELqeDnKHM9CUxlgRq6E568MGygmqqn4zr+OPvupLdYybp2PT3vz6Ewrk93
PPgLz8DBR0neYHDgk652NbVWN7JsmuajPCfSQ4m8uj9SIRPN4/M9dS3wWjAr8ilz
6338k8SlQaxG9bMV+BaSY2kQCePKF5eyIlRgejW8MRdkqSfmGg/CyY7dCz8fEzyP
/v4ZZp1CfrUjTcSrpMCxI8a6KNj45eFtcRb006nPUBAYH2JuSXVAZCXQhHarxixJ
S9ibMTkWgXr1shMoqyqOcQ5dRMy0si7uSRw6LTrtw+5+P35ESQf0fSlCul+T+z2T
ZdC93z6mwIhsUiGP4XrcpiIfSDNOiF5KkPoIspKnc1KXm4MgFlKnAuNhcQu0ugns
BKXRvF2Nk7WHrRzSY70PnktrtR9mnwYC3bJCnQ3hV0UzpZrLcSVXE+Qu63HhmGPa
QejGB3tdQDU/Uhvl0hK6CTIju/exaGErvMMNuYsZBZPdZCwjkIlbK6Ya9J8w5y3e
pjxL0T03t5GvsdcVjTkFlhMaZlp2hAAqj/4XJRkH71SZA7FGhVXbsbSmuxk9rRb2
XiDdieHq6XUv16ng/Ui6NIWxttJA12YlftESmS8218Zjco+3njkGqxnR2z4smbuy
NzNQCVRW6aGItnV4m8qK0iCdtKWOmR/6eUj/fppKsQG7GPP2Y4WqmtDbJMxJ/po7
tLM7PymibWhSqIgsF0xcQhyrOlH+jKXd6LCQ1qPDLn7tYG6iVPYF2zWa0FdzuZ7R
1m2GAG2DvcRBLqsJhpey/WMQFZYFxLcGMOvJdpBV6QW5bcxyE0rpdIrOug7qb7hT
xGYJvLoR5aELyxwHHdcfCmfsqXXthOBFbXJPvVV8adbglisiRerwP1QPYYRzhzh5
YCr8ST22vPgeVf7dtQmFOPLcft8S01+TpQl6IfAKZqebGDIU5zl+OfSOtPr0FD1f
C8CDHAyZ79nzTujqzKvxClSw4iIeT+3fyNoLwG6UFyOzHyKfE3CskxV+lVFMBjSJ
yFlU0EQFJtoncLH2vx2CRaBIi1ZGcDM6DxMQITwZDzyxYsSVQA16JsxFTovndF8g
OIMGFroEPox8nn0QYAS7f+udxytznWlDyk/cJiRoJj3aZ1TN9Mpj5HmmQ5/Y3Aja
T3zxgf1BTKxO40ycJRJfiltJQC3nmpcPm+8VlUkSaHG9GZmnNvVLB49L2zDWrM32
55OVq9sdFHrEcKWj8KOcxGDsYs67J3YTwVcbvi2jpNvkaU11OQIWiN6CRO2uJRwf
tZFAoW0mI3ZbZgD8IeW99bKO7BXKXbJh0n/hTohWJuGcKK0G9+8E5swSHSyoBFCC
v82sPeZVnZp4SkhuCyXD4m//TelzYX+/rIhY3EYXaF39obeU36ku9I3IOyK/vF8Z
+7Zu3CZrO+3/ndIEOOVpFv0cv/LgX3ttbNpoaMJZvG0ya3EuNAHcbs89xkqM0DGC
u7bUJxYQWfUhRUvllrxe8Wftdeveu/IsBrLPaeLgpYhANXU3XK+X5JK8G4OJxYTg
s2SJqVfz0xWq/0LVChQUikh3VJ+edQLMnji/LMlIOjmXhLemynNHXj4oyj12rPfS
pjEGRsWNBWaQSKXMZz5SGNtDQFt5lBthE8UUgndH1oHzsqfPA07tFLtO/cPJEcvK
Lw0yHZDBH9Ky4MhLrd8Opt/RHa8BmpLpw35GraAMelK3+itgvGqSTXciH0WyDUuI
hyIYUuT1Y7llRzYs+S/fvNNyRkeewKgz30Gg/1F8hYgGq1FuAuXAXPAFbZASwhRc
eNPLlPVW33ILbA5RUVMMCsRaJvqD1fJ0Kp3Co21VXKU9NEAY0wO4v1w74uo+v6r9
LRdXTbI9h0zUeSl252trYnm6C2wO3b+ivQXl19jA9E+xWFmtRcmFSYRLke7jB1e8
cfXxTckO7QtYXkIv8kk37LBnaGLchPc2OLvF9kiXnbE8j6HDmgPRVpvyQdSB5xCz
lw8kw21iBYTDudv999HzpBn/upihbDhuPk/wT/qwLr7ib8ZtSRXErNvxwc/kUScz
bEEDrFdAez+l3OFbXt9a+fxAkPV+JVlXD6V4fi7AkBC8oE1+Zsny4/HvlOFuXLfH
CQuFX+R8b5Jd0zNxAh5wUuVABsORK/iG6RIfQQ/RKSjBvrWEGTXQUoAB/QzGJrb2
ue9zafp9GR6skREZfKJK9m8nWFW1BrgLLdWbSu5ccmU=
`pragma protect end_protected
