-- bus_test.vhd

-- Generated using ACDS version 21.1 842

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity bus_test is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity bus_test;

architecture rtl of bus_test is
	component simple_SDC_sm is
		generic (
			DATA_WIDTH : integer := 8;
			ADDR_WIDTH : integer := 7
		);
		port (
			clk                                 : in  std_logic                    := 'X';             -- clk
			avs_s0_address                      : in  std_logic_vector(7 downto 0) := (others => 'X'); -- address
			avs_s0_waitrequest                  : out std_logic;                                       -- waitrequest
			avs_s0_read_target_synapse_addr     : in  std_logic                    := 'X';             -- read
			avs_s0_readdata_target_synapse_addr : out std_logic_vector(7 downto 0);                    -- readdata
			rst                                 : in  std_logic                    := 'X'              -- reset
		);
	end component simple_SDC_sm;

	component simple_up_server_sm is
		generic (
			DATA_WIDTH : integer := 8;
			ADDR_WIDTH : integer := 7
		);
		port (
			clk                                 : in  std_logic                    := 'X';             -- clk
			avs_s0_address                      : in  std_logic_vector(7 downto 0) := (others => 'X'); -- address
			avs_s0_write_spike                  : in  std_logic                    := 'X';             -- write
			avs_s0_writedata_spike_time         : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			avm_m0_address                      : out std_logic_vector(7 downto 0);                    -- address
			avm_m0_waitrequest                  : in  std_logic                    := 'X';             -- waitrequest
			avm_m0_write_spike                  : out std_logic;                                       -- write
			avm_m0_writedata_spike_time         : out std_logic_vector(8 downto 0);                    -- writedata
			avm_m1_address                      : out std_logic_vector(7 downto 0);                    -- address
			avm_m1_waitrequest                  : in  std_logic                    := 'X';             -- waitrequest
			avm_m1_read_target_synapse_addr     : out std_logic;                                       -- read
			avm_m1_readdata_target_synapse_addr : in  std_logic_vector(7 downto 0) := (others => 'X'); -- readdata
			rst                                 : in  std_logic                    := 'X'              -- reset
		);
	end component simple_up_server_sm;

	component simple_soma_sm is
		generic (
			THRESHOLD             : integer                      := 10;
			DATA_WIDTH            : integer                      := 8;
			ADDR_WIDTH            : integer                      := 7;
			UPLOAD_SERVER_ADDRESS : std_logic_vector(7 downto 0) := "00000001"
		);
		port (
			clk                         : in  std_logic                    := 'X';             -- clk
			avs_s0_address              : in  std_logic_vector(7 downto 0) := (others => 'X'); -- address
			avs_s0_write_synapse        : in  std_logic                    := 'X';             -- write
			avs_s0_writedata_synapse    : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			rst                         : in  std_logic                    := 'X';             -- reset
			avm_m0_address              : out std_logic_vector(7 downto 0);                    -- address
			avm_m0_waitrequest          : in  std_logic                    := 'X';             -- waitrequest
			avm_m0_write_spike          : out std_logic;                                       -- write
			avm_m0_writedata_spike_time : out std_logic_vector(7 downto 0)                     -- writedata
		);
	end component simple_soma_sm;

	component bus_test_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                           : in  std_logic                    := 'X';             -- clk
			simple_soma_SM_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                    := 'X';             -- reset
			simple_soma_SM_0_m0_address                             : in  std_logic_vector(7 downto 0) := (others => 'X'); -- address
			simple_soma_SM_0_m0_waitrequest                         : out std_logic;                                       -- waitrequest
			simple_soma_SM_0_m0_write                               : in  std_logic                    := 'X';             -- write
			simple_soma_SM_0_m0_writedata                           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			simple_UP_Server_State_Machine_0_s0_address             : out std_logic_vector(7 downto 0);                    -- address
			simple_UP_Server_State_Machine_0_s0_write               : out std_logic;                                       -- write
			simple_UP_Server_State_Machine_0_s0_writedata           : out std_logic_vector(7 downto 0)                     -- writedata
		);
	end component bus_test_mm_interconnect_0;

	component bus_test_mm_interconnect_1 is
		port (
			clk_0_clk_clk                                                           : in  std_logic                    := 'X';             -- clk
			simple_UP_Server_State_Machine_0_reset_sink_reset_bridge_in_reset_reset : in  std_logic                    := 'X';             -- reset
			simple_UP_Server_State_Machine_0_m1_address                             : in  std_logic_vector(7 downto 0) := (others => 'X'); -- address
			simple_UP_Server_State_Machine_0_m1_waitrequest                         : out std_logic;                                       -- waitrequest
			simple_UP_Server_State_Machine_0_m1_read                                : in  std_logic                    := 'X';             -- read
			simple_UP_Server_State_Machine_0_m1_readdata                            : out std_logic_vector(7 downto 0);                    -- readdata
			simple_SDC_State_Machine_0_s0_address                                   : out std_logic_vector(7 downto 0);                    -- address
			simple_SDC_State_Machine_0_s0_read                                      : out std_logic;                                       -- read
			simple_SDC_State_Machine_0_s0_readdata                                  : in  std_logic_vector(7 downto 0) := (others => 'X'); -- readdata
			simple_SDC_State_Machine_0_s0_waitrequest                               : in  std_logic                    := 'X'              -- waitrequest
		);
	end component bus_test_mm_interconnect_1;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal simple_soma_sm_0_m0_waitrequest                                 : std_logic;                    -- mm_interconnect_0:simple_soma_SM_0_m0_waitrequest -> simple_soma_SM_0:avm_m0_waitrequest
	signal simple_soma_sm_0_m0_address                                     : std_logic_vector(7 downto 0); -- simple_soma_SM_0:avm_m0_address -> mm_interconnect_0:simple_soma_SM_0_m0_address
	signal simple_soma_sm_0_m0_write                                       : std_logic;                    -- simple_soma_SM_0:avm_m0_write_spike -> mm_interconnect_0:simple_soma_SM_0_m0_write
	signal simple_soma_sm_0_m0_writedata                                   : std_logic_vector(7 downto 0); -- simple_soma_SM_0:avm_m0_writedata_spike_time -> mm_interconnect_0:simple_soma_SM_0_m0_writedata
	signal mm_interconnect_0_simple_up_server_state_machine_0_s0_address   : std_logic_vector(7 downto 0); -- mm_interconnect_0:simple_UP_Server_State_Machine_0_s0_address -> simple_UP_Server_State_Machine_0:avs_s0_address
	signal mm_interconnect_0_simple_up_server_state_machine_0_s0_write     : std_logic;                    -- mm_interconnect_0:simple_UP_Server_State_Machine_0_s0_write -> simple_UP_Server_State_Machine_0:avs_s0_write_spike
	signal mm_interconnect_0_simple_up_server_state_machine_0_s0_writedata : std_logic_vector(7 downto 0); -- mm_interconnect_0:simple_UP_Server_State_Machine_0_s0_writedata -> simple_UP_Server_State_Machine_0:avs_s0_writedata_spike_time
	signal simple_up_server_state_machine_0_m1_waitrequest                 : std_logic;                    -- mm_interconnect_1:simple_UP_Server_State_Machine_0_m1_waitrequest -> simple_UP_Server_State_Machine_0:avm_m1_waitrequest
	signal simple_up_server_state_machine_0_m1_readdata                    : std_logic_vector(7 downto 0); -- mm_interconnect_1:simple_UP_Server_State_Machine_0_m1_readdata -> simple_UP_Server_State_Machine_0:avm_m1_readdata_target_synapse_addr
	signal simple_up_server_state_machine_0_m1_address                     : std_logic_vector(7 downto 0); -- simple_UP_Server_State_Machine_0:avm_m1_address -> mm_interconnect_1:simple_UP_Server_State_Machine_0_m1_address
	signal simple_up_server_state_machine_0_m1_read                        : std_logic;                    -- simple_UP_Server_State_Machine_0:avm_m1_read_target_synapse_addr -> mm_interconnect_1:simple_UP_Server_State_Machine_0_m1_read
	signal mm_interconnect_1_simple_sdc_state_machine_0_s0_readdata        : std_logic_vector(7 downto 0); -- simple_SDC_State_Machine_0:avs_s0_readdata_target_synapse_addr -> mm_interconnect_1:simple_SDC_State_Machine_0_s0_readdata
	signal mm_interconnect_1_simple_sdc_state_machine_0_s0_waitrequest     : std_logic;                    -- simple_SDC_State_Machine_0:avs_s0_waitrequest -> mm_interconnect_1:simple_SDC_State_Machine_0_s0_waitrequest
	signal mm_interconnect_1_simple_sdc_state_machine_0_s0_address         : std_logic_vector(7 downto 0); -- mm_interconnect_1:simple_SDC_State_Machine_0_s0_address -> simple_SDC_State_Machine_0:avs_s0_address
	signal mm_interconnect_1_simple_sdc_state_machine_0_s0_read            : std_logic;                    -- mm_interconnect_1:simple_SDC_State_Machine_0_s0_read -> simple_SDC_State_Machine_0:avs_s0_read_target_synapse_addr
	signal rst_controller_reset_out_reset                                  : std_logic;                    -- rst_controller:reset_out -> [mm_interconnect_0:simple_soma_SM_0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:simple_UP_Server_State_Machine_0_reset_sink_reset_bridge_in_reset_reset, simple_SDC_State_Machine_0:rst, simple_UP_Server_State_Machine_0:rst, simple_soma_SM_0:rst]
	signal reset_reset_n_ports_inv                                         : std_logic;                    -- reset_reset_n:inv -> rst_controller:reset_in0

begin

	simple_sdc_state_machine_0 : component simple_SDC_sm
		generic map (
			DATA_WIDTH => 8,
			ADDR_WIDTH => 7
		)
		port map (
			clk                                 => clk_clk,                                                     --      clock.clk
			avs_s0_address                      => mm_interconnect_1_simple_sdc_state_machine_0_s0_address,     --         s0.address
			avs_s0_waitrequest                  => mm_interconnect_1_simple_sdc_state_machine_0_s0_waitrequest, --           .waitrequest
			avs_s0_read_target_synapse_addr     => mm_interconnect_1_simple_sdc_state_machine_0_s0_read,        --           .read
			avs_s0_readdata_target_synapse_addr => mm_interconnect_1_simple_sdc_state_machine_0_s0_readdata,    --           .readdata
			rst                                 => rst_controller_reset_out_reset                               -- reset_sink.reset
		);

	simple_up_server_state_machine_0 : component simple_up_server_sm
		generic map (
			DATA_WIDTH => 8,
			ADDR_WIDTH => 7
		)
		port map (
			clk                                 => clk_clk,                                                         --      clock.clk
			avs_s0_address                      => mm_interconnect_0_simple_up_server_state_machine_0_s0_address,   --         s0.address
			avs_s0_write_spike                  => mm_interconnect_0_simple_up_server_state_machine_0_s0_write,     --           .write
			avs_s0_writedata_spike_time         => mm_interconnect_0_simple_up_server_state_machine_0_s0_writedata, --           .writedata
			avm_m0_address                      => open,                                                            --         m0.address
			avm_m0_waitrequest                  => open,                                                            --           .waitrequest
			avm_m0_write_spike                  => open,                                                            --           .write
			avm_m0_writedata_spike_time         => open,                                                            --           .writedata
			avm_m1_address                      => simple_up_server_state_machine_0_m1_address,                     --         m1.address
			avm_m1_waitrequest                  => simple_up_server_state_machine_0_m1_waitrequest,                 --           .waitrequest
			avm_m1_read_target_synapse_addr     => simple_up_server_state_machine_0_m1_read,                        --           .read
			avm_m1_readdata_target_synapse_addr => simple_up_server_state_machine_0_m1_readdata,                    --           .readdata
			rst                                 => rst_controller_reset_out_reset                                   -- reset_sink.reset
		);

	simple_soma_sm_0 : component simple_soma_sm
		generic map (
			THRESHOLD             => 10,
			DATA_WIDTH            => 8,
			ADDR_WIDTH            => 7,
			UPLOAD_SERVER_ADDRESS => "00000001"
		)
		port map (
			clk                         => clk_clk,                         --      clock.clk
			avs_s0_address              => open,                            --         s0.address
			avs_s0_write_synapse        => open,                            --           .write
			avs_s0_writedata_synapse    => open,                            --           .writedata
			rst                         => rst_controller_reset_out_reset,  -- reset_sink.reset
			avm_m0_address              => simple_soma_sm_0_m0_address,     --         m0.address
			avm_m0_waitrequest          => simple_soma_sm_0_m0_waitrequest, --           .waitrequest
			avm_m0_write_spike          => simple_soma_sm_0_m0_write,       --           .write
			avm_m0_writedata_spike_time => simple_soma_sm_0_m0_writedata    --           .writedata
		);

	mm_interconnect_0 : component bus_test_mm_interconnect_0
		port map (
			clk_0_clk_clk                                           => clk_clk,                                                         --                                         clk_0_clk.clk
			simple_soma_SM_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                  -- simple_soma_SM_0_reset_sink_reset_bridge_in_reset.reset
			simple_soma_SM_0_m0_address                             => simple_soma_sm_0_m0_address,                                     --                               simple_soma_SM_0_m0.address
			simple_soma_SM_0_m0_waitrequest                         => simple_soma_sm_0_m0_waitrequest,                                 --                                                  .waitrequest
			simple_soma_SM_0_m0_write                               => simple_soma_sm_0_m0_write,                                       --                                                  .write
			simple_soma_SM_0_m0_writedata                           => simple_soma_sm_0_m0_writedata,                                   --                                                  .writedata
			simple_UP_Server_State_Machine_0_s0_address             => mm_interconnect_0_simple_up_server_state_machine_0_s0_address,   --               simple_UP_Server_State_Machine_0_s0.address
			simple_UP_Server_State_Machine_0_s0_write               => mm_interconnect_0_simple_up_server_state_machine_0_s0_write,     --                                                  .write
			simple_UP_Server_State_Machine_0_s0_writedata           => mm_interconnect_0_simple_up_server_state_machine_0_s0_writedata  --                                                  .writedata
		);

	mm_interconnect_1 : component bus_test_mm_interconnect_1
		port map (
			clk_0_clk_clk                                                           => clk_clk,                                                     --                                                         clk_0_clk.clk
			simple_UP_Server_State_Machine_0_reset_sink_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                              -- simple_UP_Server_State_Machine_0_reset_sink_reset_bridge_in_reset.reset
			simple_UP_Server_State_Machine_0_m1_address                             => simple_up_server_state_machine_0_m1_address,                 --                               simple_UP_Server_State_Machine_0_m1.address
			simple_UP_Server_State_Machine_0_m1_waitrequest                         => simple_up_server_state_machine_0_m1_waitrequest,             --                                                                  .waitrequest
			simple_UP_Server_State_Machine_0_m1_read                                => simple_up_server_state_machine_0_m1_read,                    --                                                                  .read
			simple_UP_Server_State_Machine_0_m1_readdata                            => simple_up_server_state_machine_0_m1_readdata,                --                                                                  .readdata
			simple_SDC_State_Machine_0_s0_address                                   => mm_interconnect_1_simple_sdc_state_machine_0_s0_address,     --                                     simple_SDC_State_Machine_0_s0.address
			simple_SDC_State_Machine_0_s0_read                                      => mm_interconnect_1_simple_sdc_state_machine_0_s0_read,        --                                                                  .read
			simple_SDC_State_Machine_0_s0_readdata                                  => mm_interconnect_1_simple_sdc_state_machine_0_s0_readdata,    --                                                                  .readdata
			simple_SDC_State_Machine_0_s0_waitrequest                               => mm_interconnect_1_simple_sdc_state_machine_0_s0_waitrequest  --                                                                  .waitrequest
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

end architecture rtl; -- of bus_test
